library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.math_real.all;
use work.constants_pkg.ALL;

package lut_pkg is
    constant SINE_FS : LUT := (
   0 => to_unsigned(512, AMPLITUDE_WIDTH),
   1 => to_unsigned(512, AMPLITUDE_WIDTH),
   2 => to_unsigned(513, AMPLITUDE_WIDTH),
   3 => to_unsigned(514, AMPLITUDE_WIDTH),
   4 => to_unsigned(515, AMPLITUDE_WIDTH),
   5 => to_unsigned(515, AMPLITUDE_WIDTH),
   6 => to_unsigned(516, AMPLITUDE_WIDTH),
   7 => to_unsigned(517, AMPLITUDE_WIDTH),
   8 => to_unsigned(518, AMPLITUDE_WIDTH),
   9 => to_unsigned(519, AMPLITUDE_WIDTH),
  10 => to_unsigned(519, AMPLITUDE_WIDTH),
  11 => to_unsigned(520, AMPLITUDE_WIDTH),
  12 => to_unsigned(521, AMPLITUDE_WIDTH),
  13 => to_unsigned(522, AMPLITUDE_WIDTH),
  14 => to_unsigned(522, AMPLITUDE_WIDTH),
  15 => to_unsigned(523, AMPLITUDE_WIDTH),
  16 => to_unsigned(524, AMPLITUDE_WIDTH),
  17 => to_unsigned(525, AMPLITUDE_WIDTH),
  18 => to_unsigned(526, AMPLITUDE_WIDTH),
  19 => to_unsigned(526, AMPLITUDE_WIDTH),
  20 => to_unsigned(527, AMPLITUDE_WIDTH),
  21 => to_unsigned(528, AMPLITUDE_WIDTH),
  22 => to_unsigned(529, AMPLITUDE_WIDTH),
  23 => to_unsigned(530, AMPLITUDE_WIDTH),
  24 => to_unsigned(530, AMPLITUDE_WIDTH),
  25 => to_unsigned(531, AMPLITUDE_WIDTH),
  26 => to_unsigned(532, AMPLITUDE_WIDTH),
  27 => to_unsigned(533, AMPLITUDE_WIDTH),
  28 => to_unsigned(533, AMPLITUDE_WIDTH),
  29 => to_unsigned(534, AMPLITUDE_WIDTH),
  30 => to_unsigned(535, AMPLITUDE_WIDTH),
  31 => to_unsigned(536, AMPLITUDE_WIDTH),
  32 => to_unsigned(537, AMPLITUDE_WIDTH),
  33 => to_unsigned(537, AMPLITUDE_WIDTH),
  34 => to_unsigned(538, AMPLITUDE_WIDTH),
  35 => to_unsigned(539, AMPLITUDE_WIDTH),
  36 => to_unsigned(540, AMPLITUDE_WIDTH),
  37 => to_unsigned(541, AMPLITUDE_WIDTH),
  38 => to_unsigned(541, AMPLITUDE_WIDTH),
  39 => to_unsigned(542, AMPLITUDE_WIDTH),
  40 => to_unsigned(543, AMPLITUDE_WIDTH),
  41 => to_unsigned(544, AMPLITUDE_WIDTH),
  42 => to_unsigned(544, AMPLITUDE_WIDTH),
  43 => to_unsigned(545, AMPLITUDE_WIDTH),
  44 => to_unsigned(546, AMPLITUDE_WIDTH),
  45 => to_unsigned(547, AMPLITUDE_WIDTH),
  46 => to_unsigned(548, AMPLITUDE_WIDTH),
  47 => to_unsigned(548, AMPLITUDE_WIDTH),
  48 => to_unsigned(549, AMPLITUDE_WIDTH),
  49 => to_unsigned(550, AMPLITUDE_WIDTH),
  50 => to_unsigned(551, AMPLITUDE_WIDTH),
  51 => to_unsigned(552, AMPLITUDE_WIDTH),
  52 => to_unsigned(552, AMPLITUDE_WIDTH),
  53 => to_unsigned(553, AMPLITUDE_WIDTH),
  54 => to_unsigned(554, AMPLITUDE_WIDTH),
  55 => to_unsigned(555, AMPLITUDE_WIDTH),
  56 => to_unsigned(555, AMPLITUDE_WIDTH),
  57 => to_unsigned(556, AMPLITUDE_WIDTH),
  58 => to_unsigned(557, AMPLITUDE_WIDTH),
  59 => to_unsigned(558, AMPLITUDE_WIDTH),
  60 => to_unsigned(559, AMPLITUDE_WIDTH),
  61 => to_unsigned(559, AMPLITUDE_WIDTH),
  62 => to_unsigned(560, AMPLITUDE_WIDTH),
  63 => to_unsigned(561, AMPLITUDE_WIDTH),
  64 => to_unsigned(562, AMPLITUDE_WIDTH),
  65 => to_unsigned(562, AMPLITUDE_WIDTH),
  66 => to_unsigned(563, AMPLITUDE_WIDTH),
  67 => to_unsigned(564, AMPLITUDE_WIDTH),
  68 => to_unsigned(565, AMPLITUDE_WIDTH),
  69 => to_unsigned(566, AMPLITUDE_WIDTH),
  70 => to_unsigned(566, AMPLITUDE_WIDTH),
  71 => to_unsigned(567, AMPLITUDE_WIDTH),
  72 => to_unsigned(568, AMPLITUDE_WIDTH),
  73 => to_unsigned(569, AMPLITUDE_WIDTH),
  74 => to_unsigned(569, AMPLITUDE_WIDTH),
  75 => to_unsigned(570, AMPLITUDE_WIDTH),
  76 => to_unsigned(571, AMPLITUDE_WIDTH),
  77 => to_unsigned(572, AMPLITUDE_WIDTH),
  78 => to_unsigned(573, AMPLITUDE_WIDTH),
  79 => to_unsigned(573, AMPLITUDE_WIDTH),
  80 => to_unsigned(574, AMPLITUDE_WIDTH),
  81 => to_unsigned(575, AMPLITUDE_WIDTH),
  82 => to_unsigned(576, AMPLITUDE_WIDTH),
  83 => to_unsigned(577, AMPLITUDE_WIDTH),
  84 => to_unsigned(577, AMPLITUDE_WIDTH),
  85 => to_unsigned(578, AMPLITUDE_WIDTH),
  86 => to_unsigned(579, AMPLITUDE_WIDTH),
  87 => to_unsigned(580, AMPLITUDE_WIDTH),
  88 => to_unsigned(580, AMPLITUDE_WIDTH),
  89 => to_unsigned(581, AMPLITUDE_WIDTH),
  90 => to_unsigned(582, AMPLITUDE_WIDTH),
  91 => to_unsigned(583, AMPLITUDE_WIDTH),
  92 => to_unsigned(584, AMPLITUDE_WIDTH),
  93 => to_unsigned(584, AMPLITUDE_WIDTH),
  94 => to_unsigned(585, AMPLITUDE_WIDTH),
  95 => to_unsigned(586, AMPLITUDE_WIDTH),
  96 => to_unsigned(587, AMPLITUDE_WIDTH),
  97 => to_unsigned(587, AMPLITUDE_WIDTH),
  98 => to_unsigned(588, AMPLITUDE_WIDTH),
  99 => to_unsigned(589, AMPLITUDE_WIDTH),
 100 => to_unsigned(590, AMPLITUDE_WIDTH),
 101 => to_unsigned(591, AMPLITUDE_WIDTH),
 102 => to_unsigned(591, AMPLITUDE_WIDTH),
 103 => to_unsigned(592, AMPLITUDE_WIDTH),
 104 => to_unsigned(593, AMPLITUDE_WIDTH),
 105 => to_unsigned(594, AMPLITUDE_WIDTH),
 106 => to_unsigned(594, AMPLITUDE_WIDTH),
 107 => to_unsigned(595, AMPLITUDE_WIDTH),
 108 => to_unsigned(596, AMPLITUDE_WIDTH),
 109 => to_unsigned(597, AMPLITUDE_WIDTH),
 110 => to_unsigned(597, AMPLITUDE_WIDTH),
 111 => to_unsigned(598, AMPLITUDE_WIDTH),
 112 => to_unsigned(599, AMPLITUDE_WIDTH),
 113 => to_unsigned(600, AMPLITUDE_WIDTH),
 114 => to_unsigned(601, AMPLITUDE_WIDTH),
 115 => to_unsigned(601, AMPLITUDE_WIDTH),
 116 => to_unsigned(602, AMPLITUDE_WIDTH),
 117 => to_unsigned(603, AMPLITUDE_WIDTH),
 118 => to_unsigned(604, AMPLITUDE_WIDTH),
 119 => to_unsigned(604, AMPLITUDE_WIDTH),
 120 => to_unsigned(605, AMPLITUDE_WIDTH),
 121 => to_unsigned(606, AMPLITUDE_WIDTH),
 122 => to_unsigned(607, AMPLITUDE_WIDTH),
 123 => to_unsigned(608, AMPLITUDE_WIDTH),
 124 => to_unsigned(608, AMPLITUDE_WIDTH),
 125 => to_unsigned(609, AMPLITUDE_WIDTH),
 126 => to_unsigned(610, AMPLITUDE_WIDTH),
 127 => to_unsigned(611, AMPLITUDE_WIDTH),
 128 => to_unsigned(611, AMPLITUDE_WIDTH),
 129 => to_unsigned(612, AMPLITUDE_WIDTH),
 130 => to_unsigned(613, AMPLITUDE_WIDTH),
 131 => to_unsigned(614, AMPLITUDE_WIDTH),
 132 => to_unsigned(614, AMPLITUDE_WIDTH),
 133 => to_unsigned(615, AMPLITUDE_WIDTH),
 134 => to_unsigned(616, AMPLITUDE_WIDTH),
 135 => to_unsigned(617, AMPLITUDE_WIDTH),
 136 => to_unsigned(618, AMPLITUDE_WIDTH),
 137 => to_unsigned(618, AMPLITUDE_WIDTH),
 138 => to_unsigned(619, AMPLITUDE_WIDTH),
 139 => to_unsigned(620, AMPLITUDE_WIDTH),
 140 => to_unsigned(621, AMPLITUDE_WIDTH),
 141 => to_unsigned(621, AMPLITUDE_WIDTH),
 142 => to_unsigned(622, AMPLITUDE_WIDTH),
 143 => to_unsigned(623, AMPLITUDE_WIDTH),
 144 => to_unsigned(624, AMPLITUDE_WIDTH),
 145 => to_unsigned(624, AMPLITUDE_WIDTH),
 146 => to_unsigned(625, AMPLITUDE_WIDTH),
 147 => to_unsigned(626, AMPLITUDE_WIDTH),
 148 => to_unsigned(627, AMPLITUDE_WIDTH),
 149 => to_unsigned(628, AMPLITUDE_WIDTH),
 150 => to_unsigned(628, AMPLITUDE_WIDTH),
 151 => to_unsigned(629, AMPLITUDE_WIDTH),
 152 => to_unsigned(630, AMPLITUDE_WIDTH),
 153 => to_unsigned(631, AMPLITUDE_WIDTH),
 154 => to_unsigned(631, AMPLITUDE_WIDTH),
 155 => to_unsigned(632, AMPLITUDE_WIDTH),
 156 => to_unsigned(633, AMPLITUDE_WIDTH),
 157 => to_unsigned(634, AMPLITUDE_WIDTH),
 158 => to_unsigned(634, AMPLITUDE_WIDTH),
 159 => to_unsigned(635, AMPLITUDE_WIDTH),
 160 => to_unsigned(636, AMPLITUDE_WIDTH),
 161 => to_unsigned(637, AMPLITUDE_WIDTH),
 162 => to_unsigned(637, AMPLITUDE_WIDTH),
 163 => to_unsigned(638, AMPLITUDE_WIDTH),
 164 => to_unsigned(639, AMPLITUDE_WIDTH),
 165 => to_unsigned(640, AMPLITUDE_WIDTH),
 166 => to_unsigned(640, AMPLITUDE_WIDTH),
 167 => to_unsigned(641, AMPLITUDE_WIDTH),
 168 => to_unsigned(642, AMPLITUDE_WIDTH),
 169 => to_unsigned(643, AMPLITUDE_WIDTH),
 170 => to_unsigned(644, AMPLITUDE_WIDTH),
 171 => to_unsigned(644, AMPLITUDE_WIDTH),
 172 => to_unsigned(645, AMPLITUDE_WIDTH),
 173 => to_unsigned(646, AMPLITUDE_WIDTH),
 174 => to_unsigned(647, AMPLITUDE_WIDTH),
 175 => to_unsigned(647, AMPLITUDE_WIDTH),
 176 => to_unsigned(648, AMPLITUDE_WIDTH),
 177 => to_unsigned(649, AMPLITUDE_WIDTH),
 178 => to_unsigned(650, AMPLITUDE_WIDTH),
 179 => to_unsigned(650, AMPLITUDE_WIDTH),
 180 => to_unsigned(651, AMPLITUDE_WIDTH),
 181 => to_unsigned(652, AMPLITUDE_WIDTH),
 182 => to_unsigned(653, AMPLITUDE_WIDTH),
 183 => to_unsigned(653, AMPLITUDE_WIDTH),
 184 => to_unsigned(654, AMPLITUDE_WIDTH),
 185 => to_unsigned(655, AMPLITUDE_WIDTH),
 186 => to_unsigned(656, AMPLITUDE_WIDTH),
 187 => to_unsigned(656, AMPLITUDE_WIDTH),
 188 => to_unsigned(657, AMPLITUDE_WIDTH),
 189 => to_unsigned(658, AMPLITUDE_WIDTH),
 190 => to_unsigned(659, AMPLITUDE_WIDTH),
 191 => to_unsigned(659, AMPLITUDE_WIDTH),
 192 => to_unsigned(660, AMPLITUDE_WIDTH),
 193 => to_unsigned(661, AMPLITUDE_WIDTH),
 194 => to_unsigned(662, AMPLITUDE_WIDTH),
 195 => to_unsigned(662, AMPLITUDE_WIDTH),
 196 => to_unsigned(663, AMPLITUDE_WIDTH),
 197 => to_unsigned(664, AMPLITUDE_WIDTH),
 198 => to_unsigned(665, AMPLITUDE_WIDTH),
 199 => to_unsigned(665, AMPLITUDE_WIDTH),
 200 => to_unsigned(666, AMPLITUDE_WIDTH),
 201 => to_unsigned(667, AMPLITUDE_WIDTH),
 202 => to_unsigned(668, AMPLITUDE_WIDTH),
 203 => to_unsigned(668, AMPLITUDE_WIDTH),
 204 => to_unsigned(669, AMPLITUDE_WIDTH),
 205 => to_unsigned(670, AMPLITUDE_WIDTH),
 206 => to_unsigned(671, AMPLITUDE_WIDTH),
 207 => to_unsigned(671, AMPLITUDE_WIDTH),
 208 => to_unsigned(672, AMPLITUDE_WIDTH),
 209 => to_unsigned(673, AMPLITUDE_WIDTH),
 210 => to_unsigned(674, AMPLITUDE_WIDTH),
 211 => to_unsigned(674, AMPLITUDE_WIDTH),
 212 => to_unsigned(675, AMPLITUDE_WIDTH),
 213 => to_unsigned(676, AMPLITUDE_WIDTH),
 214 => to_unsigned(677, AMPLITUDE_WIDTH),
 215 => to_unsigned(677, AMPLITUDE_WIDTH),
 216 => to_unsigned(678, AMPLITUDE_WIDTH),
 217 => to_unsigned(679, AMPLITUDE_WIDTH),
 218 => to_unsigned(680, AMPLITUDE_WIDTH),
 219 => to_unsigned(680, AMPLITUDE_WIDTH),
 220 => to_unsigned(681, AMPLITUDE_WIDTH),
 221 => to_unsigned(682, AMPLITUDE_WIDTH),
 222 => to_unsigned(683, AMPLITUDE_WIDTH),
 223 => to_unsigned(683, AMPLITUDE_WIDTH),
 224 => to_unsigned(684, AMPLITUDE_WIDTH),
 225 => to_unsigned(685, AMPLITUDE_WIDTH),
 226 => to_unsigned(685, AMPLITUDE_WIDTH),
 227 => to_unsigned(686, AMPLITUDE_WIDTH),
 228 => to_unsigned(687, AMPLITUDE_WIDTH),
 229 => to_unsigned(688, AMPLITUDE_WIDTH),
 230 => to_unsigned(688, AMPLITUDE_WIDTH),
 231 => to_unsigned(689, AMPLITUDE_WIDTH),
 232 => to_unsigned(690, AMPLITUDE_WIDTH),
 233 => to_unsigned(691, AMPLITUDE_WIDTH),
 234 => to_unsigned(691, AMPLITUDE_WIDTH),
 235 => to_unsigned(692, AMPLITUDE_WIDTH),
 236 => to_unsigned(693, AMPLITUDE_WIDTH),
 237 => to_unsigned(694, AMPLITUDE_WIDTH),
 238 => to_unsigned(694, AMPLITUDE_WIDTH),
 239 => to_unsigned(695, AMPLITUDE_WIDTH),
 240 => to_unsigned(696, AMPLITUDE_WIDTH),
 241 => to_unsigned(696, AMPLITUDE_WIDTH),
 242 => to_unsigned(697, AMPLITUDE_WIDTH),
 243 => to_unsigned(698, AMPLITUDE_WIDTH),
 244 => to_unsigned(699, AMPLITUDE_WIDTH),
 245 => to_unsigned(699, AMPLITUDE_WIDTH),
 246 => to_unsigned(700, AMPLITUDE_WIDTH),
 247 => to_unsigned(701, AMPLITUDE_WIDTH),
 248 => to_unsigned(702, AMPLITUDE_WIDTH),
 249 => to_unsigned(702, AMPLITUDE_WIDTH),
 250 => to_unsigned(703, AMPLITUDE_WIDTH),
 251 => to_unsigned(704, AMPLITUDE_WIDTH),
 252 => to_unsigned(705, AMPLITUDE_WIDTH),
 253 => to_unsigned(705, AMPLITUDE_WIDTH),
 254 => to_unsigned(706, AMPLITUDE_WIDTH),
 255 => to_unsigned(707, AMPLITUDE_WIDTH),
 256 => to_unsigned(707, AMPLITUDE_WIDTH),
 257 => to_unsigned(708, AMPLITUDE_WIDTH),
 258 => to_unsigned(709, AMPLITUDE_WIDTH),
 259 => to_unsigned(710, AMPLITUDE_WIDTH),
 260 => to_unsigned(710, AMPLITUDE_WIDTH),
 261 => to_unsigned(711, AMPLITUDE_WIDTH),
 262 => to_unsigned(712, AMPLITUDE_WIDTH),
 263 => to_unsigned(712, AMPLITUDE_WIDTH),
 264 => to_unsigned(713, AMPLITUDE_WIDTH),
 265 => to_unsigned(714, AMPLITUDE_WIDTH),
 266 => to_unsigned(715, AMPLITUDE_WIDTH),
 267 => to_unsigned(715, AMPLITUDE_WIDTH),
 268 => to_unsigned(716, AMPLITUDE_WIDTH),
 269 => to_unsigned(717, AMPLITUDE_WIDTH),
 270 => to_unsigned(718, AMPLITUDE_WIDTH),
 271 => to_unsigned(718, AMPLITUDE_WIDTH),
 272 => to_unsigned(719, AMPLITUDE_WIDTH),
 273 => to_unsigned(720, AMPLITUDE_WIDTH),
 274 => to_unsigned(720, AMPLITUDE_WIDTH),
 275 => to_unsigned(721, AMPLITUDE_WIDTH),
 276 => to_unsigned(722, AMPLITUDE_WIDTH),
 277 => to_unsigned(723, AMPLITUDE_WIDTH),
 278 => to_unsigned(723, AMPLITUDE_WIDTH),
 279 => to_unsigned(724, AMPLITUDE_WIDTH),
 280 => to_unsigned(725, AMPLITUDE_WIDTH),
 281 => to_unsigned(725, AMPLITUDE_WIDTH),
 282 => to_unsigned(726, AMPLITUDE_WIDTH),
 283 => to_unsigned(727, AMPLITUDE_WIDTH),
 284 => to_unsigned(728, AMPLITUDE_WIDTH),
 285 => to_unsigned(728, AMPLITUDE_WIDTH),
 286 => to_unsigned(729, AMPLITUDE_WIDTH),
 287 => to_unsigned(730, AMPLITUDE_WIDTH),
 288 => to_unsigned(730, AMPLITUDE_WIDTH),
 289 => to_unsigned(731, AMPLITUDE_WIDTH),
 290 => to_unsigned(732, AMPLITUDE_WIDTH),
 291 => to_unsigned(733, AMPLITUDE_WIDTH),
 292 => to_unsigned(733, AMPLITUDE_WIDTH),
 293 => to_unsigned(734, AMPLITUDE_WIDTH),
 294 => to_unsigned(735, AMPLITUDE_WIDTH),
 295 => to_unsigned(735, AMPLITUDE_WIDTH),
 296 => to_unsigned(736, AMPLITUDE_WIDTH),
 297 => to_unsigned(737, AMPLITUDE_WIDTH),
 298 => to_unsigned(737, AMPLITUDE_WIDTH),
 299 => to_unsigned(738, AMPLITUDE_WIDTH),
 300 => to_unsigned(739, AMPLITUDE_WIDTH),
 301 => to_unsigned(740, AMPLITUDE_WIDTH),
 302 => to_unsigned(740, AMPLITUDE_WIDTH),
 303 => to_unsigned(741, AMPLITUDE_WIDTH),
 304 => to_unsigned(742, AMPLITUDE_WIDTH),
 305 => to_unsigned(742, AMPLITUDE_WIDTH),
 306 => to_unsigned(743, AMPLITUDE_WIDTH),
 307 => to_unsigned(744, AMPLITUDE_WIDTH),
 308 => to_unsigned(744, AMPLITUDE_WIDTH),
 309 => to_unsigned(745, AMPLITUDE_WIDTH),
 310 => to_unsigned(746, AMPLITUDE_WIDTH),
 311 => to_unsigned(747, AMPLITUDE_WIDTH),
 312 => to_unsigned(747, AMPLITUDE_WIDTH),
 313 => to_unsigned(748, AMPLITUDE_WIDTH),
 314 => to_unsigned(749, AMPLITUDE_WIDTH),
 315 => to_unsigned(749, AMPLITUDE_WIDTH),
 316 => to_unsigned(750, AMPLITUDE_WIDTH),
 317 => to_unsigned(751, AMPLITUDE_WIDTH),
 318 => to_unsigned(751, AMPLITUDE_WIDTH),
 319 => to_unsigned(752, AMPLITUDE_WIDTH),
 320 => to_unsigned(753, AMPLITUDE_WIDTH),
 321 => to_unsigned(754, AMPLITUDE_WIDTH),
 322 => to_unsigned(754, AMPLITUDE_WIDTH),
 323 => to_unsigned(755, AMPLITUDE_WIDTH),
 324 => to_unsigned(756, AMPLITUDE_WIDTH),
 325 => to_unsigned(756, AMPLITUDE_WIDTH),
 326 => to_unsigned(757, AMPLITUDE_WIDTH),
 327 => to_unsigned(758, AMPLITUDE_WIDTH),
 328 => to_unsigned(758, AMPLITUDE_WIDTH),
 329 => to_unsigned(759, AMPLITUDE_WIDTH),
 330 => to_unsigned(760, AMPLITUDE_WIDTH),
 331 => to_unsigned(760, AMPLITUDE_WIDTH),
 332 => to_unsigned(761, AMPLITUDE_WIDTH),
 333 => to_unsigned(762, AMPLITUDE_WIDTH),
 334 => to_unsigned(762, AMPLITUDE_WIDTH),
 335 => to_unsigned(763, AMPLITUDE_WIDTH),
 336 => to_unsigned(764, AMPLITUDE_WIDTH),
 337 => to_unsigned(765, AMPLITUDE_WIDTH),
 338 => to_unsigned(765, AMPLITUDE_WIDTH),
 339 => to_unsigned(766, AMPLITUDE_WIDTH),
 340 => to_unsigned(767, AMPLITUDE_WIDTH),
 341 => to_unsigned(767, AMPLITUDE_WIDTH),
 342 => to_unsigned(768, AMPLITUDE_WIDTH),
 343 => to_unsigned(769, AMPLITUDE_WIDTH),
 344 => to_unsigned(769, AMPLITUDE_WIDTH),
 345 => to_unsigned(770, AMPLITUDE_WIDTH),
 346 => to_unsigned(771, AMPLITUDE_WIDTH),
 347 => to_unsigned(771, AMPLITUDE_WIDTH),
 348 => to_unsigned(772, AMPLITUDE_WIDTH),
 349 => to_unsigned(773, AMPLITUDE_WIDTH),
 350 => to_unsigned(773, AMPLITUDE_WIDTH),
 351 => to_unsigned(774, AMPLITUDE_WIDTH),
 352 => to_unsigned(775, AMPLITUDE_WIDTH),
 353 => to_unsigned(775, AMPLITUDE_WIDTH),
 354 => to_unsigned(776, AMPLITUDE_WIDTH),
 355 => to_unsigned(777, AMPLITUDE_WIDTH),
 356 => to_unsigned(777, AMPLITUDE_WIDTH),
 357 => to_unsigned(778, AMPLITUDE_WIDTH),
 358 => to_unsigned(779, AMPLITUDE_WIDTH),
 359 => to_unsigned(779, AMPLITUDE_WIDTH),
 360 => to_unsigned(780, AMPLITUDE_WIDTH),
 361 => to_unsigned(781, AMPLITUDE_WIDTH),
 362 => to_unsigned(781, AMPLITUDE_WIDTH),
 363 => to_unsigned(782, AMPLITUDE_WIDTH),
 364 => to_unsigned(783, AMPLITUDE_WIDTH),
 365 => to_unsigned(783, AMPLITUDE_WIDTH),
 366 => to_unsigned(784, AMPLITUDE_WIDTH),
 367 => to_unsigned(785, AMPLITUDE_WIDTH),
 368 => to_unsigned(785, AMPLITUDE_WIDTH),
 369 => to_unsigned(786, AMPLITUDE_WIDTH),
 370 => to_unsigned(787, AMPLITUDE_WIDTH),
 371 => to_unsigned(787, AMPLITUDE_WIDTH),
 372 => to_unsigned(788, AMPLITUDE_WIDTH),
 373 => to_unsigned(789, AMPLITUDE_WIDTH),
 374 => to_unsigned(789, AMPLITUDE_WIDTH),
 375 => to_unsigned(790, AMPLITUDE_WIDTH),
 376 => to_unsigned(791, AMPLITUDE_WIDTH),
 377 => to_unsigned(791, AMPLITUDE_WIDTH),
 378 => to_unsigned(792, AMPLITUDE_WIDTH),
 379 => to_unsigned(793, AMPLITUDE_WIDTH),
 380 => to_unsigned(793, AMPLITUDE_WIDTH),
 381 => to_unsigned(794, AMPLITUDE_WIDTH),
 382 => to_unsigned(795, AMPLITUDE_WIDTH),
 383 => to_unsigned(795, AMPLITUDE_WIDTH),
 384 => to_unsigned(796, AMPLITUDE_WIDTH),
 385 => to_unsigned(797, AMPLITUDE_WIDTH),
 386 => to_unsigned(797, AMPLITUDE_WIDTH),
 387 => to_unsigned(798, AMPLITUDE_WIDTH),
 388 => to_unsigned(799, AMPLITUDE_WIDTH),
 389 => to_unsigned(799, AMPLITUDE_WIDTH),
 390 => to_unsigned(800, AMPLITUDE_WIDTH),
 391 => to_unsigned(800, AMPLITUDE_WIDTH),
 392 => to_unsigned(801, AMPLITUDE_WIDTH),
 393 => to_unsigned(802, AMPLITUDE_WIDTH),
 394 => to_unsigned(802, AMPLITUDE_WIDTH),
 395 => to_unsigned(803, AMPLITUDE_WIDTH),
 396 => to_unsigned(804, AMPLITUDE_WIDTH),
 397 => to_unsigned(804, AMPLITUDE_WIDTH),
 398 => to_unsigned(805, AMPLITUDE_WIDTH),
 399 => to_unsigned(806, AMPLITUDE_WIDTH),
 400 => to_unsigned(806, AMPLITUDE_WIDTH),
 401 => to_unsigned(807, AMPLITUDE_WIDTH),
 402 => to_unsigned(808, AMPLITUDE_WIDTH),
 403 => to_unsigned(808, AMPLITUDE_WIDTH),
 404 => to_unsigned(809, AMPLITUDE_WIDTH),
 405 => to_unsigned(809, AMPLITUDE_WIDTH),
 406 => to_unsigned(810, AMPLITUDE_WIDTH),
 407 => to_unsigned(811, AMPLITUDE_WIDTH),
 408 => to_unsigned(811, AMPLITUDE_WIDTH),
 409 => to_unsigned(812, AMPLITUDE_WIDTH),
 410 => to_unsigned(813, AMPLITUDE_WIDTH),
 411 => to_unsigned(813, AMPLITUDE_WIDTH),
 412 => to_unsigned(814, AMPLITUDE_WIDTH),
 413 => to_unsigned(815, AMPLITUDE_WIDTH),
 414 => to_unsigned(815, AMPLITUDE_WIDTH),
 415 => to_unsigned(816, AMPLITUDE_WIDTH),
 416 => to_unsigned(816, AMPLITUDE_WIDTH),
 417 => to_unsigned(817, AMPLITUDE_WIDTH),
 418 => to_unsigned(818, AMPLITUDE_WIDTH),
 419 => to_unsigned(818, AMPLITUDE_WIDTH),
 420 => to_unsigned(819, AMPLITUDE_WIDTH),
 421 => to_unsigned(820, AMPLITUDE_WIDTH),
 422 => to_unsigned(820, AMPLITUDE_WIDTH),
 423 => to_unsigned(821, AMPLITUDE_WIDTH),
 424 => to_unsigned(821, AMPLITUDE_WIDTH),
 425 => to_unsigned(822, AMPLITUDE_WIDTH),
 426 => to_unsigned(823, AMPLITUDE_WIDTH),
 427 => to_unsigned(823, AMPLITUDE_WIDTH),
 428 => to_unsigned(824, AMPLITUDE_WIDTH),
 429 => to_unsigned(825, AMPLITUDE_WIDTH),
 430 => to_unsigned(825, AMPLITUDE_WIDTH),
 431 => to_unsigned(826, AMPLITUDE_WIDTH),
 432 => to_unsigned(826, AMPLITUDE_WIDTH),
 433 => to_unsigned(827, AMPLITUDE_WIDTH),
 434 => to_unsigned(828, AMPLITUDE_WIDTH),
 435 => to_unsigned(828, AMPLITUDE_WIDTH),
 436 => to_unsigned(829, AMPLITUDE_WIDTH),
 437 => to_unsigned(830, AMPLITUDE_WIDTH),
 438 => to_unsigned(830, AMPLITUDE_WIDTH),
 439 => to_unsigned(831, AMPLITUDE_WIDTH),
 440 => to_unsigned(831, AMPLITUDE_WIDTH),
 441 => to_unsigned(832, AMPLITUDE_WIDTH),
 442 => to_unsigned(833, AMPLITUDE_WIDTH),
 443 => to_unsigned(833, AMPLITUDE_WIDTH),
 444 => to_unsigned(834, AMPLITUDE_WIDTH),
 445 => to_unsigned(834, AMPLITUDE_WIDTH),
 446 => to_unsigned(835, AMPLITUDE_WIDTH),
 447 => to_unsigned(836, AMPLITUDE_WIDTH),
 448 => to_unsigned(836, AMPLITUDE_WIDTH),
 449 => to_unsigned(837, AMPLITUDE_WIDTH),
 450 => to_unsigned(837, AMPLITUDE_WIDTH),
 451 => to_unsigned(838, AMPLITUDE_WIDTH),
 452 => to_unsigned(839, AMPLITUDE_WIDTH),
 453 => to_unsigned(839, AMPLITUDE_WIDTH),
 454 => to_unsigned(840, AMPLITUDE_WIDTH),
 455 => to_unsigned(840, AMPLITUDE_WIDTH),
 456 => to_unsigned(841, AMPLITUDE_WIDTH),
 457 => to_unsigned(842, AMPLITUDE_WIDTH),
 458 => to_unsigned(842, AMPLITUDE_WIDTH),
 459 => to_unsigned(843, AMPLITUDE_WIDTH),
 460 => to_unsigned(843, AMPLITUDE_WIDTH),
 461 => to_unsigned(844, AMPLITUDE_WIDTH),
 462 => to_unsigned(845, AMPLITUDE_WIDTH),
 463 => to_unsigned(845, AMPLITUDE_WIDTH),
 464 => to_unsigned(846, AMPLITUDE_WIDTH),
 465 => to_unsigned(846, AMPLITUDE_WIDTH),
 466 => to_unsigned(847, AMPLITUDE_WIDTH),
 467 => to_unsigned(848, AMPLITUDE_WIDTH),
 468 => to_unsigned(848, AMPLITUDE_WIDTH),
 469 => to_unsigned(849, AMPLITUDE_WIDTH),
 470 => to_unsigned(849, AMPLITUDE_WIDTH),
 471 => to_unsigned(850, AMPLITUDE_WIDTH),
 472 => to_unsigned(851, AMPLITUDE_WIDTH),
 473 => to_unsigned(851, AMPLITUDE_WIDTH),
 474 => to_unsigned(852, AMPLITUDE_WIDTH),
 475 => to_unsigned(852, AMPLITUDE_WIDTH),
 476 => to_unsigned(853, AMPLITUDE_WIDTH),
 477 => to_unsigned(854, AMPLITUDE_WIDTH),
 478 => to_unsigned(854, AMPLITUDE_WIDTH),
 479 => to_unsigned(855, AMPLITUDE_WIDTH),
 480 => to_unsigned(855, AMPLITUDE_WIDTH),
 481 => to_unsigned(856, AMPLITUDE_WIDTH),
 482 => to_unsigned(856, AMPLITUDE_WIDTH),
 483 => to_unsigned(857, AMPLITUDE_WIDTH),
 484 => to_unsigned(858, AMPLITUDE_WIDTH),
 485 => to_unsigned(858, AMPLITUDE_WIDTH),
 486 => to_unsigned(859, AMPLITUDE_WIDTH),
 487 => to_unsigned(859, AMPLITUDE_WIDTH),
 488 => to_unsigned(860, AMPLITUDE_WIDTH),
 489 => to_unsigned(860, AMPLITUDE_WIDTH),
 490 => to_unsigned(861, AMPLITUDE_WIDTH),
 491 => to_unsigned(862, AMPLITUDE_WIDTH),
 492 => to_unsigned(862, AMPLITUDE_WIDTH),
 493 => to_unsigned(863, AMPLITUDE_WIDTH),
 494 => to_unsigned(863, AMPLITUDE_WIDTH),
 495 => to_unsigned(864, AMPLITUDE_WIDTH),
 496 => to_unsigned(864, AMPLITUDE_WIDTH),
 497 => to_unsigned(865, AMPLITUDE_WIDTH),
 498 => to_unsigned(866, AMPLITUDE_WIDTH),
 499 => to_unsigned(866, AMPLITUDE_WIDTH),
 500 => to_unsigned(867, AMPLITUDE_WIDTH),
 501 => to_unsigned(867, AMPLITUDE_WIDTH),
 502 => to_unsigned(868, AMPLITUDE_WIDTH),
 503 => to_unsigned(868, AMPLITUDE_WIDTH),
 504 => to_unsigned(869, AMPLITUDE_WIDTH),
 505 => to_unsigned(870, AMPLITUDE_WIDTH),
 506 => to_unsigned(870, AMPLITUDE_WIDTH),
 507 => to_unsigned(871, AMPLITUDE_WIDTH),
 508 => to_unsigned(871, AMPLITUDE_WIDTH),
 509 => to_unsigned(872, AMPLITUDE_WIDTH),
 510 => to_unsigned(872, AMPLITUDE_WIDTH),
 511 => to_unsigned(873, AMPLITUDE_WIDTH),
 512 => to_unsigned(873, AMPLITUDE_WIDTH),
 513 => to_unsigned(874, AMPLITUDE_WIDTH),
 514 => to_unsigned(875, AMPLITUDE_WIDTH),
 515 => to_unsigned(875, AMPLITUDE_WIDTH),
 516 => to_unsigned(876, AMPLITUDE_WIDTH),
 517 => to_unsigned(876, AMPLITUDE_WIDTH),
 518 => to_unsigned(877, AMPLITUDE_WIDTH),
 519 => to_unsigned(877, AMPLITUDE_WIDTH),
 520 => to_unsigned(878, AMPLITUDE_WIDTH),
 521 => to_unsigned(878, AMPLITUDE_WIDTH),
 522 => to_unsigned(879, AMPLITUDE_WIDTH),
 523 => to_unsigned(880, AMPLITUDE_WIDTH),
 524 => to_unsigned(880, AMPLITUDE_WIDTH),
 525 => to_unsigned(881, AMPLITUDE_WIDTH),
 526 => to_unsigned(881, AMPLITUDE_WIDTH),
 527 => to_unsigned(882, AMPLITUDE_WIDTH),
 528 => to_unsigned(882, AMPLITUDE_WIDTH),
 529 => to_unsigned(883, AMPLITUDE_WIDTH),
 530 => to_unsigned(883, AMPLITUDE_WIDTH),
 531 => to_unsigned(884, AMPLITUDE_WIDTH),
 532 => to_unsigned(884, AMPLITUDE_WIDTH),
 533 => to_unsigned(885, AMPLITUDE_WIDTH),
 534 => to_unsigned(885, AMPLITUDE_WIDTH),
 535 => to_unsigned(886, AMPLITUDE_WIDTH),
 536 => to_unsigned(887, AMPLITUDE_WIDTH),
 537 => to_unsigned(887, AMPLITUDE_WIDTH),
 538 => to_unsigned(888, AMPLITUDE_WIDTH),
 539 => to_unsigned(888, AMPLITUDE_WIDTH),
 540 => to_unsigned(889, AMPLITUDE_WIDTH),
 541 => to_unsigned(889, AMPLITUDE_WIDTH),
 542 => to_unsigned(890, AMPLITUDE_WIDTH),
 543 => to_unsigned(890, AMPLITUDE_WIDTH),
 544 => to_unsigned(891, AMPLITUDE_WIDTH),
 545 => to_unsigned(891, AMPLITUDE_WIDTH),
 546 => to_unsigned(892, AMPLITUDE_WIDTH),
 547 => to_unsigned(892, AMPLITUDE_WIDTH),
 548 => to_unsigned(893, AMPLITUDE_WIDTH),
 549 => to_unsigned(893, AMPLITUDE_WIDTH),
 550 => to_unsigned(894, AMPLITUDE_WIDTH),
 551 => to_unsigned(894, AMPLITUDE_WIDTH),
 552 => to_unsigned(895, AMPLITUDE_WIDTH),
 553 => to_unsigned(895, AMPLITUDE_WIDTH),
 554 => to_unsigned(896, AMPLITUDE_WIDTH),
 555 => to_unsigned(897, AMPLITUDE_WIDTH),
 556 => to_unsigned(897, AMPLITUDE_WIDTH),
 557 => to_unsigned(898, AMPLITUDE_WIDTH),
 558 => to_unsigned(898, AMPLITUDE_WIDTH),
 559 => to_unsigned(899, AMPLITUDE_WIDTH),
 560 => to_unsigned(899, AMPLITUDE_WIDTH),
 561 => to_unsigned(900, AMPLITUDE_WIDTH),
 562 => to_unsigned(900, AMPLITUDE_WIDTH),
 563 => to_unsigned(901, AMPLITUDE_WIDTH),
 564 => to_unsigned(901, AMPLITUDE_WIDTH),
 565 => to_unsigned(902, AMPLITUDE_WIDTH),
 566 => to_unsigned(902, AMPLITUDE_WIDTH),
 567 => to_unsigned(903, AMPLITUDE_WIDTH),
 568 => to_unsigned(903, AMPLITUDE_WIDTH),
 569 => to_unsigned(904, AMPLITUDE_WIDTH),
 570 => to_unsigned(904, AMPLITUDE_WIDTH),
 571 => to_unsigned(905, AMPLITUDE_WIDTH),
 572 => to_unsigned(905, AMPLITUDE_WIDTH),
 573 => to_unsigned(906, AMPLITUDE_WIDTH),
 574 => to_unsigned(906, AMPLITUDE_WIDTH),
 575 => to_unsigned(907, AMPLITUDE_WIDTH),
 576 => to_unsigned(907, AMPLITUDE_WIDTH),
 577 => to_unsigned(908, AMPLITUDE_WIDTH),
 578 => to_unsigned(908, AMPLITUDE_WIDTH),
 579 => to_unsigned(909, AMPLITUDE_WIDTH),
 580 => to_unsigned(909, AMPLITUDE_WIDTH),
 581 => to_unsigned(910, AMPLITUDE_WIDTH),
 582 => to_unsigned(910, AMPLITUDE_WIDTH),
 583 => to_unsigned(911, AMPLITUDE_WIDTH),
 584 => to_unsigned(911, AMPLITUDE_WIDTH),
 585 => to_unsigned(912, AMPLITUDE_WIDTH),
 586 => to_unsigned(912, AMPLITUDE_WIDTH),
 587 => to_unsigned(913, AMPLITUDE_WIDTH),
 588 => to_unsigned(913, AMPLITUDE_WIDTH),
 589 => to_unsigned(914, AMPLITUDE_WIDTH),
 590 => to_unsigned(914, AMPLITUDE_WIDTH),
 591 => to_unsigned(915, AMPLITUDE_WIDTH),
 592 => to_unsigned(915, AMPLITUDE_WIDTH),
 593 => to_unsigned(916, AMPLITUDE_WIDTH),
 594 => to_unsigned(916, AMPLITUDE_WIDTH),
 595 => to_unsigned(916, AMPLITUDE_WIDTH),
 596 => to_unsigned(917, AMPLITUDE_WIDTH),
 597 => to_unsigned(917, AMPLITUDE_WIDTH),
 598 => to_unsigned(918, AMPLITUDE_WIDTH),
 599 => to_unsigned(918, AMPLITUDE_WIDTH),
 600 => to_unsigned(919, AMPLITUDE_WIDTH),
 601 => to_unsigned(919, AMPLITUDE_WIDTH),
 602 => to_unsigned(920, AMPLITUDE_WIDTH),
 603 => to_unsigned(920, AMPLITUDE_WIDTH),
 604 => to_unsigned(921, AMPLITUDE_WIDTH),
 605 => to_unsigned(921, AMPLITUDE_WIDTH),
 606 => to_unsigned(922, AMPLITUDE_WIDTH),
 607 => to_unsigned(922, AMPLITUDE_WIDTH),
 608 => to_unsigned(923, AMPLITUDE_WIDTH),
 609 => to_unsigned(923, AMPLITUDE_WIDTH),
 610 => to_unsigned(924, AMPLITUDE_WIDTH),
 611 => to_unsigned(924, AMPLITUDE_WIDTH),
 612 => to_unsigned(924, AMPLITUDE_WIDTH),
 613 => to_unsigned(925, AMPLITUDE_WIDTH),
 614 => to_unsigned(925, AMPLITUDE_WIDTH),
 615 => to_unsigned(926, AMPLITUDE_WIDTH),
 616 => to_unsigned(926, AMPLITUDE_WIDTH),
 617 => to_unsigned(927, AMPLITUDE_WIDTH),
 618 => to_unsigned(927, AMPLITUDE_WIDTH),
 619 => to_unsigned(928, AMPLITUDE_WIDTH),
 620 => to_unsigned(928, AMPLITUDE_WIDTH),
 621 => to_unsigned(929, AMPLITUDE_WIDTH),
 622 => to_unsigned(929, AMPLITUDE_WIDTH),
 623 => to_unsigned(930, AMPLITUDE_WIDTH),
 624 => to_unsigned(930, AMPLITUDE_WIDTH),
 625 => to_unsigned(930, AMPLITUDE_WIDTH),
 626 => to_unsigned(931, AMPLITUDE_WIDTH),
 627 => to_unsigned(931, AMPLITUDE_WIDTH),
 628 => to_unsigned(932, AMPLITUDE_WIDTH),
 629 => to_unsigned(932, AMPLITUDE_WIDTH),
 630 => to_unsigned(933, AMPLITUDE_WIDTH),
 631 => to_unsigned(933, AMPLITUDE_WIDTH),
 632 => to_unsigned(934, AMPLITUDE_WIDTH),
 633 => to_unsigned(934, AMPLITUDE_WIDTH),
 634 => to_unsigned(934, AMPLITUDE_WIDTH),
 635 => to_unsigned(935, AMPLITUDE_WIDTH),
 636 => to_unsigned(935, AMPLITUDE_WIDTH),
 637 => to_unsigned(936, AMPLITUDE_WIDTH),
 638 => to_unsigned(936, AMPLITUDE_WIDTH),
 639 => to_unsigned(937, AMPLITUDE_WIDTH),
 640 => to_unsigned(937, AMPLITUDE_WIDTH),
 641 => to_unsigned(938, AMPLITUDE_WIDTH),
 642 => to_unsigned(938, AMPLITUDE_WIDTH),
 643 => to_unsigned(938, AMPLITUDE_WIDTH),
 644 => to_unsigned(939, AMPLITUDE_WIDTH),
 645 => to_unsigned(939, AMPLITUDE_WIDTH),
 646 => to_unsigned(940, AMPLITUDE_WIDTH),
 647 => to_unsigned(940, AMPLITUDE_WIDTH),
 648 => to_unsigned(941, AMPLITUDE_WIDTH),
 649 => to_unsigned(941, AMPLITUDE_WIDTH),
 650 => to_unsigned(941, AMPLITUDE_WIDTH),
 651 => to_unsigned(942, AMPLITUDE_WIDTH),
 652 => to_unsigned(942, AMPLITUDE_WIDTH),
 653 => to_unsigned(943, AMPLITUDE_WIDTH),
 654 => to_unsigned(943, AMPLITUDE_WIDTH),
 655 => to_unsigned(943, AMPLITUDE_WIDTH),
 656 => to_unsigned(944, AMPLITUDE_WIDTH),
 657 => to_unsigned(944, AMPLITUDE_WIDTH),
 658 => to_unsigned(945, AMPLITUDE_WIDTH),
 659 => to_unsigned(945, AMPLITUDE_WIDTH),
 660 => to_unsigned(946, AMPLITUDE_WIDTH),
 661 => to_unsigned(946, AMPLITUDE_WIDTH),
 662 => to_unsigned(946, AMPLITUDE_WIDTH),
 663 => to_unsigned(947, AMPLITUDE_WIDTH),
 664 => to_unsigned(947, AMPLITUDE_WIDTH),
 665 => to_unsigned(948, AMPLITUDE_WIDTH),
 666 => to_unsigned(948, AMPLITUDE_WIDTH),
 667 => to_unsigned(948, AMPLITUDE_WIDTH),
 668 => to_unsigned(949, AMPLITUDE_WIDTH),
 669 => to_unsigned(949, AMPLITUDE_WIDTH),
 670 => to_unsigned(950, AMPLITUDE_WIDTH),
 671 => to_unsigned(950, AMPLITUDE_WIDTH),
 672 => to_unsigned(950, AMPLITUDE_WIDTH),
 673 => to_unsigned(951, AMPLITUDE_WIDTH),
 674 => to_unsigned(951, AMPLITUDE_WIDTH),
 675 => to_unsigned(952, AMPLITUDE_WIDTH),
 676 => to_unsigned(952, AMPLITUDE_WIDTH),
 677 => to_unsigned(952, AMPLITUDE_WIDTH),
 678 => to_unsigned(953, AMPLITUDE_WIDTH),
 679 => to_unsigned(953, AMPLITUDE_WIDTH),
 680 => to_unsigned(954, AMPLITUDE_WIDTH),
 681 => to_unsigned(954, AMPLITUDE_WIDTH),
 682 => to_unsigned(954, AMPLITUDE_WIDTH),
 683 => to_unsigned(955, AMPLITUDE_WIDTH),
 684 => to_unsigned(955, AMPLITUDE_WIDTH),
 685 => to_unsigned(956, AMPLITUDE_WIDTH),
 686 => to_unsigned(956, AMPLITUDE_WIDTH),
 687 => to_unsigned(956, AMPLITUDE_WIDTH),
 688 => to_unsigned(957, AMPLITUDE_WIDTH),
 689 => to_unsigned(957, AMPLITUDE_WIDTH),
 690 => to_unsigned(958, AMPLITUDE_WIDTH),
 691 => to_unsigned(958, AMPLITUDE_WIDTH),
 692 => to_unsigned(958, AMPLITUDE_WIDTH),
 693 => to_unsigned(959, AMPLITUDE_WIDTH),
 694 => to_unsigned(959, AMPLITUDE_WIDTH),
 695 => to_unsigned(959, AMPLITUDE_WIDTH),
 696 => to_unsigned(960, AMPLITUDE_WIDTH),
 697 => to_unsigned(960, AMPLITUDE_WIDTH),
 698 => to_unsigned(961, AMPLITUDE_WIDTH),
 699 => to_unsigned(961, AMPLITUDE_WIDTH),
 700 => to_unsigned(961, AMPLITUDE_WIDTH),
 701 => to_unsigned(962, AMPLITUDE_WIDTH),
 702 => to_unsigned(962, AMPLITUDE_WIDTH),
 703 => to_unsigned(962, AMPLITUDE_WIDTH),
 704 => to_unsigned(963, AMPLITUDE_WIDTH),
 705 => to_unsigned(963, AMPLITUDE_WIDTH),
 706 => to_unsigned(964, AMPLITUDE_WIDTH),
 707 => to_unsigned(964, AMPLITUDE_WIDTH),
 708 => to_unsigned(964, AMPLITUDE_WIDTH),
 709 => to_unsigned(965, AMPLITUDE_WIDTH),
 710 => to_unsigned(965, AMPLITUDE_WIDTH),
 711 => to_unsigned(965, AMPLITUDE_WIDTH),
 712 => to_unsigned(966, AMPLITUDE_WIDTH),
 713 => to_unsigned(966, AMPLITUDE_WIDTH),
 714 => to_unsigned(966, AMPLITUDE_WIDTH),
 715 => to_unsigned(967, AMPLITUDE_WIDTH),
 716 => to_unsigned(967, AMPLITUDE_WIDTH),
 717 => to_unsigned(968, AMPLITUDE_WIDTH),
 718 => to_unsigned(968, AMPLITUDE_WIDTH),
 719 => to_unsigned(968, AMPLITUDE_WIDTH),
 720 => to_unsigned(969, AMPLITUDE_WIDTH),
 721 => to_unsigned(969, AMPLITUDE_WIDTH),
 722 => to_unsigned(969, AMPLITUDE_WIDTH),
 723 => to_unsigned(970, AMPLITUDE_WIDTH),
 724 => to_unsigned(970, AMPLITUDE_WIDTH),
 725 => to_unsigned(970, AMPLITUDE_WIDTH),
 726 => to_unsigned(971, AMPLITUDE_WIDTH),
 727 => to_unsigned(971, AMPLITUDE_WIDTH),
 728 => to_unsigned(971, AMPLITUDE_WIDTH),
 729 => to_unsigned(972, AMPLITUDE_WIDTH),
 730 => to_unsigned(972, AMPLITUDE_WIDTH),
 731 => to_unsigned(972, AMPLITUDE_WIDTH),
 732 => to_unsigned(973, AMPLITUDE_WIDTH),
 733 => to_unsigned(973, AMPLITUDE_WIDTH),
 734 => to_unsigned(973, AMPLITUDE_WIDTH),
 735 => to_unsigned(974, AMPLITUDE_WIDTH),
 736 => to_unsigned(974, AMPLITUDE_WIDTH),
 737 => to_unsigned(974, AMPLITUDE_WIDTH),
 738 => to_unsigned(975, AMPLITUDE_WIDTH),
 739 => to_unsigned(975, AMPLITUDE_WIDTH),
 740 => to_unsigned(975, AMPLITUDE_WIDTH),
 741 => to_unsigned(976, AMPLITUDE_WIDTH),
 742 => to_unsigned(976, AMPLITUDE_WIDTH),
 743 => to_unsigned(976, AMPLITUDE_WIDTH),
 744 => to_unsigned(977, AMPLITUDE_WIDTH),
 745 => to_unsigned(977, AMPLITUDE_WIDTH),
 746 => to_unsigned(977, AMPLITUDE_WIDTH),
 747 => to_unsigned(978, AMPLITUDE_WIDTH),
 748 => to_unsigned(978, AMPLITUDE_WIDTH),
 749 => to_unsigned(978, AMPLITUDE_WIDTH),
 750 => to_unsigned(979, AMPLITUDE_WIDTH),
 751 => to_unsigned(979, AMPLITUDE_WIDTH),
 752 => to_unsigned(979, AMPLITUDE_WIDTH),
 753 => to_unsigned(980, AMPLITUDE_WIDTH),
 754 => to_unsigned(980, AMPLITUDE_WIDTH),
 755 => to_unsigned(980, AMPLITUDE_WIDTH),
 756 => to_unsigned(981, AMPLITUDE_WIDTH),
 757 => to_unsigned(981, AMPLITUDE_WIDTH),
 758 => to_unsigned(981, AMPLITUDE_WIDTH),
 759 => to_unsigned(982, AMPLITUDE_WIDTH),
 760 => to_unsigned(982, AMPLITUDE_WIDTH),
 761 => to_unsigned(982, AMPLITUDE_WIDTH),
 762 => to_unsigned(982, AMPLITUDE_WIDTH),
 763 => to_unsigned(983, AMPLITUDE_WIDTH),
 764 => to_unsigned(983, AMPLITUDE_WIDTH),
 765 => to_unsigned(983, AMPLITUDE_WIDTH),
 766 => to_unsigned(984, AMPLITUDE_WIDTH),
 767 => to_unsigned(984, AMPLITUDE_WIDTH),
 768 => to_unsigned(984, AMPLITUDE_WIDTH),
 769 => to_unsigned(985, AMPLITUDE_WIDTH),
 770 => to_unsigned(985, AMPLITUDE_WIDTH),
 771 => to_unsigned(985, AMPLITUDE_WIDTH),
 772 => to_unsigned(985, AMPLITUDE_WIDTH),
 773 => to_unsigned(986, AMPLITUDE_WIDTH),
 774 => to_unsigned(986, AMPLITUDE_WIDTH),
 775 => to_unsigned(986, AMPLITUDE_WIDTH),
 776 => to_unsigned(987, AMPLITUDE_WIDTH),
 777 => to_unsigned(987, AMPLITUDE_WIDTH),
 778 => to_unsigned(987, AMPLITUDE_WIDTH),
 779 => to_unsigned(988, AMPLITUDE_WIDTH),
 780 => to_unsigned(988, AMPLITUDE_WIDTH),
 781 => to_unsigned(988, AMPLITUDE_WIDTH),
 782 => to_unsigned(988, AMPLITUDE_WIDTH),
 783 => to_unsigned(989, AMPLITUDE_WIDTH),
 784 => to_unsigned(989, AMPLITUDE_WIDTH),
 785 => to_unsigned(989, AMPLITUDE_WIDTH),
 786 => to_unsigned(990, AMPLITUDE_WIDTH),
 787 => to_unsigned(990, AMPLITUDE_WIDTH),
 788 => to_unsigned(990, AMPLITUDE_WIDTH),
 789 => to_unsigned(990, AMPLITUDE_WIDTH),
 790 => to_unsigned(991, AMPLITUDE_WIDTH),
 791 => to_unsigned(991, AMPLITUDE_WIDTH),
 792 => to_unsigned(991, AMPLITUDE_WIDTH),
 793 => to_unsigned(991, AMPLITUDE_WIDTH),
 794 => to_unsigned(992, AMPLITUDE_WIDTH),
 795 => to_unsigned(992, AMPLITUDE_WIDTH),
 796 => to_unsigned(992, AMPLITUDE_WIDTH),
 797 => to_unsigned(993, AMPLITUDE_WIDTH),
 798 => to_unsigned(993, AMPLITUDE_WIDTH),
 799 => to_unsigned(993, AMPLITUDE_WIDTH),
 800 => to_unsigned(993, AMPLITUDE_WIDTH),
 801 => to_unsigned(994, AMPLITUDE_WIDTH),
 802 => to_unsigned(994, AMPLITUDE_WIDTH),
 803 => to_unsigned(994, AMPLITUDE_WIDTH),
 804 => to_unsigned(994, AMPLITUDE_WIDTH),
 805 => to_unsigned(995, AMPLITUDE_WIDTH),
 806 => to_unsigned(995, AMPLITUDE_WIDTH),
 807 => to_unsigned(995, AMPLITUDE_WIDTH),
 808 => to_unsigned(995, AMPLITUDE_WIDTH),
 809 => to_unsigned(996, AMPLITUDE_WIDTH),
 810 => to_unsigned(996, AMPLITUDE_WIDTH),
 811 => to_unsigned(996, AMPLITUDE_WIDTH),
 812 => to_unsigned(996, AMPLITUDE_WIDTH),
 813 => to_unsigned(997, AMPLITUDE_WIDTH),
 814 => to_unsigned(997, AMPLITUDE_WIDTH),
 815 => to_unsigned(997, AMPLITUDE_WIDTH),
 816 => to_unsigned(997, AMPLITUDE_WIDTH),
 817 => to_unsigned(998, AMPLITUDE_WIDTH),
 818 => to_unsigned(998, AMPLITUDE_WIDTH),
 819 => to_unsigned(998, AMPLITUDE_WIDTH),
 820 => to_unsigned(998, AMPLITUDE_WIDTH),
 821 => to_unsigned(999, AMPLITUDE_WIDTH),
 822 => to_unsigned(999, AMPLITUDE_WIDTH),
 823 => to_unsigned(999, AMPLITUDE_WIDTH),
 824 => to_unsigned(999, AMPLITUDE_WIDTH),
 825 => to_unsigned(1000, AMPLITUDE_WIDTH),
 826 => to_unsigned(1000, AMPLITUDE_WIDTH),
 827 => to_unsigned(1000, AMPLITUDE_WIDTH),
 828 => to_unsigned(1000, AMPLITUDE_WIDTH),
 829 => to_unsigned(1000, AMPLITUDE_WIDTH),
 830 => to_unsigned(1001, AMPLITUDE_WIDTH),
 831 => to_unsigned(1001, AMPLITUDE_WIDTH),
 832 => to_unsigned(1001, AMPLITUDE_WIDTH),
 833 => to_unsigned(1001, AMPLITUDE_WIDTH),
 834 => to_unsigned(1002, AMPLITUDE_WIDTH),
 835 => to_unsigned(1002, AMPLITUDE_WIDTH),
 836 => to_unsigned(1002, AMPLITUDE_WIDTH),
 837 => to_unsigned(1002, AMPLITUDE_WIDTH),
 838 => to_unsigned(1003, AMPLITUDE_WIDTH),
 839 => to_unsigned(1003, AMPLITUDE_WIDTH),
 840 => to_unsigned(1003, AMPLITUDE_WIDTH),
 841 => to_unsigned(1003, AMPLITUDE_WIDTH),
 842 => to_unsigned(1003, AMPLITUDE_WIDTH),
 843 => to_unsigned(1004, AMPLITUDE_WIDTH),
 844 => to_unsigned(1004, AMPLITUDE_WIDTH),
 845 => to_unsigned(1004, AMPLITUDE_WIDTH),
 846 => to_unsigned(1004, AMPLITUDE_WIDTH),
 847 => to_unsigned(1004, AMPLITUDE_WIDTH),
 848 => to_unsigned(1005, AMPLITUDE_WIDTH),
 849 => to_unsigned(1005, AMPLITUDE_WIDTH),
 850 => to_unsigned(1005, AMPLITUDE_WIDTH),
 851 => to_unsigned(1005, AMPLITUDE_WIDTH),
 852 => to_unsigned(1005, AMPLITUDE_WIDTH),
 853 => to_unsigned(1006, AMPLITUDE_WIDTH),
 854 => to_unsigned(1006, AMPLITUDE_WIDTH),
 855 => to_unsigned(1006, AMPLITUDE_WIDTH),
 856 => to_unsigned(1006, AMPLITUDE_WIDTH),
 857 => to_unsigned(1006, AMPLITUDE_WIDTH),
 858 => to_unsigned(1007, AMPLITUDE_WIDTH),
 859 => to_unsigned(1007, AMPLITUDE_WIDTH),
 860 => to_unsigned(1007, AMPLITUDE_WIDTH),
 861 => to_unsigned(1007, AMPLITUDE_WIDTH),
 862 => to_unsigned(1007, AMPLITUDE_WIDTH),
 863 => to_unsigned(1008, AMPLITUDE_WIDTH),
 864 => to_unsigned(1008, AMPLITUDE_WIDTH),
 865 => to_unsigned(1008, AMPLITUDE_WIDTH),
 866 => to_unsigned(1008, AMPLITUDE_WIDTH),
 867 => to_unsigned(1008, AMPLITUDE_WIDTH),
 868 => to_unsigned(1009, AMPLITUDE_WIDTH),
 869 => to_unsigned(1009, AMPLITUDE_WIDTH),
 870 => to_unsigned(1009, AMPLITUDE_WIDTH),
 871 => to_unsigned(1009, AMPLITUDE_WIDTH),
 872 => to_unsigned(1009, AMPLITUDE_WIDTH),
 873 => to_unsigned(1009, AMPLITUDE_WIDTH),
 874 => to_unsigned(1010, AMPLITUDE_WIDTH),
 875 => to_unsigned(1010, AMPLITUDE_WIDTH),
 876 => to_unsigned(1010, AMPLITUDE_WIDTH),
 877 => to_unsigned(1010, AMPLITUDE_WIDTH),
 878 => to_unsigned(1010, AMPLITUDE_WIDTH),
 879 => to_unsigned(1011, AMPLITUDE_WIDTH),
 880 => to_unsigned(1011, AMPLITUDE_WIDTH),
 881 => to_unsigned(1011, AMPLITUDE_WIDTH),
 882 => to_unsigned(1011, AMPLITUDE_WIDTH),
 883 => to_unsigned(1011, AMPLITUDE_WIDTH),
 884 => to_unsigned(1011, AMPLITUDE_WIDTH),
 885 => to_unsigned(1012, AMPLITUDE_WIDTH),
 886 => to_unsigned(1012, AMPLITUDE_WIDTH),
 887 => to_unsigned(1012, AMPLITUDE_WIDTH),
 888 => to_unsigned(1012, AMPLITUDE_WIDTH),
 889 => to_unsigned(1012, AMPLITUDE_WIDTH),
 890 => to_unsigned(1012, AMPLITUDE_WIDTH),
 891 => to_unsigned(1013, AMPLITUDE_WIDTH),
 892 => to_unsigned(1013, AMPLITUDE_WIDTH),
 893 => to_unsigned(1013, AMPLITUDE_WIDTH),
 894 => to_unsigned(1013, AMPLITUDE_WIDTH),
 895 => to_unsigned(1013, AMPLITUDE_WIDTH),
 896 => to_unsigned(1013, AMPLITUDE_WIDTH),
 897 => to_unsigned(1013, AMPLITUDE_WIDTH),
 898 => to_unsigned(1014, AMPLITUDE_WIDTH),
 899 => to_unsigned(1014, AMPLITUDE_WIDTH),
 900 => to_unsigned(1014, AMPLITUDE_WIDTH),
 901 => to_unsigned(1014, AMPLITUDE_WIDTH),
 902 => to_unsigned(1014, AMPLITUDE_WIDTH),
 903 => to_unsigned(1014, AMPLITUDE_WIDTH),
 904 => to_unsigned(1014, AMPLITUDE_WIDTH),
 905 => to_unsigned(1015, AMPLITUDE_WIDTH),
 906 => to_unsigned(1015, AMPLITUDE_WIDTH),
 907 => to_unsigned(1015, AMPLITUDE_WIDTH),
 908 => to_unsigned(1015, AMPLITUDE_WIDTH),
 909 => to_unsigned(1015, AMPLITUDE_WIDTH),
 910 => to_unsigned(1015, AMPLITUDE_WIDTH),
 911 => to_unsigned(1015, AMPLITUDE_WIDTH),
 912 => to_unsigned(1016, AMPLITUDE_WIDTH),
 913 => to_unsigned(1016, AMPLITUDE_WIDTH),
 914 => to_unsigned(1016, AMPLITUDE_WIDTH),
 915 => to_unsigned(1016, AMPLITUDE_WIDTH),
 916 => to_unsigned(1016, AMPLITUDE_WIDTH),
 917 => to_unsigned(1016, AMPLITUDE_WIDTH),
 918 => to_unsigned(1016, AMPLITUDE_WIDTH),
 919 => to_unsigned(1016, AMPLITUDE_WIDTH),
 920 => to_unsigned(1017, AMPLITUDE_WIDTH),
 921 => to_unsigned(1017, AMPLITUDE_WIDTH),
 922 => to_unsigned(1017, AMPLITUDE_WIDTH),
 923 => to_unsigned(1017, AMPLITUDE_WIDTH),
 924 => to_unsigned(1017, AMPLITUDE_WIDTH),
 925 => to_unsigned(1017, AMPLITUDE_WIDTH),
 926 => to_unsigned(1017, AMPLITUDE_WIDTH),
 927 => to_unsigned(1017, AMPLITUDE_WIDTH),
 928 => to_unsigned(1018, AMPLITUDE_WIDTH),
 929 => to_unsigned(1018, AMPLITUDE_WIDTH),
 930 => to_unsigned(1018, AMPLITUDE_WIDTH),
 931 => to_unsigned(1018, AMPLITUDE_WIDTH),
 932 => to_unsigned(1018, AMPLITUDE_WIDTH),
 933 => to_unsigned(1018, AMPLITUDE_WIDTH),
 934 => to_unsigned(1018, AMPLITUDE_WIDTH),
 935 => to_unsigned(1018, AMPLITUDE_WIDTH),
 936 => to_unsigned(1018, AMPLITUDE_WIDTH),
 937 => to_unsigned(1019, AMPLITUDE_WIDTH),
 938 => to_unsigned(1019, AMPLITUDE_WIDTH),
 939 => to_unsigned(1019, AMPLITUDE_WIDTH),
 940 => to_unsigned(1019, AMPLITUDE_WIDTH),
 941 => to_unsigned(1019, AMPLITUDE_WIDTH),
 942 => to_unsigned(1019, AMPLITUDE_WIDTH),
 943 => to_unsigned(1019, AMPLITUDE_WIDTH),
 944 => to_unsigned(1019, AMPLITUDE_WIDTH),
 945 => to_unsigned(1019, AMPLITUDE_WIDTH),
 946 => to_unsigned(1019, AMPLITUDE_WIDTH),
 947 => to_unsigned(1020, AMPLITUDE_WIDTH),
 948 => to_unsigned(1020, AMPLITUDE_WIDTH),
 949 => to_unsigned(1020, AMPLITUDE_WIDTH),
 950 => to_unsigned(1020, AMPLITUDE_WIDTH),
 951 => to_unsigned(1020, AMPLITUDE_WIDTH),
 952 => to_unsigned(1020, AMPLITUDE_WIDTH),
 953 => to_unsigned(1020, AMPLITUDE_WIDTH),
 954 => to_unsigned(1020, AMPLITUDE_WIDTH),
 955 => to_unsigned(1020, AMPLITUDE_WIDTH),
 956 => to_unsigned(1020, AMPLITUDE_WIDTH),
 957 => to_unsigned(1020, AMPLITUDE_WIDTH),
 958 => to_unsigned(1020, AMPLITUDE_WIDTH),
 959 => to_unsigned(1021, AMPLITUDE_WIDTH),
 960 => to_unsigned(1021, AMPLITUDE_WIDTH),
 961 => to_unsigned(1021, AMPLITUDE_WIDTH),
 962 => to_unsigned(1021, AMPLITUDE_WIDTH),
 963 => to_unsigned(1021, AMPLITUDE_WIDTH),
 964 => to_unsigned(1021, AMPLITUDE_WIDTH),
 965 => to_unsigned(1021, AMPLITUDE_WIDTH),
 966 => to_unsigned(1021, AMPLITUDE_WIDTH),
 967 => to_unsigned(1021, AMPLITUDE_WIDTH),
 968 => to_unsigned(1021, AMPLITUDE_WIDTH),
 969 => to_unsigned(1021, AMPLITUDE_WIDTH),
 970 => to_unsigned(1021, AMPLITUDE_WIDTH),
 971 => to_unsigned(1021, AMPLITUDE_WIDTH),
 972 => to_unsigned(1021, AMPLITUDE_WIDTH),
 973 => to_unsigned(1021, AMPLITUDE_WIDTH),
 974 => to_unsigned(1022, AMPLITUDE_WIDTH),
 975 => to_unsigned(1022, AMPLITUDE_WIDTH),
 976 => to_unsigned(1022, AMPLITUDE_WIDTH),
 977 => to_unsigned(1022, AMPLITUDE_WIDTH),
 978 => to_unsigned(1022, AMPLITUDE_WIDTH),
 979 => to_unsigned(1022, AMPLITUDE_WIDTH),
 980 => to_unsigned(1022, AMPLITUDE_WIDTH),
 981 => to_unsigned(1022, AMPLITUDE_WIDTH),
 982 => to_unsigned(1022, AMPLITUDE_WIDTH),
 983 => to_unsigned(1022, AMPLITUDE_WIDTH),
 984 => to_unsigned(1022, AMPLITUDE_WIDTH),
 985 => to_unsigned(1022, AMPLITUDE_WIDTH),
 986 => to_unsigned(1022, AMPLITUDE_WIDTH),
 987 => to_unsigned(1022, AMPLITUDE_WIDTH),
 988 => to_unsigned(1022, AMPLITUDE_WIDTH),
 989 => to_unsigned(1022, AMPLITUDE_WIDTH),
 990 => to_unsigned(1022, AMPLITUDE_WIDTH),
 991 => to_unsigned(1022, AMPLITUDE_WIDTH),
 992 => to_unsigned(1022, AMPLITUDE_WIDTH),
 993 => to_unsigned(1022, AMPLITUDE_WIDTH),
 994 => to_unsigned(1022, AMPLITUDE_WIDTH),
 995 => to_unsigned(1023, AMPLITUDE_WIDTH),
 996 => to_unsigned(1023, AMPLITUDE_WIDTH),
 997 => to_unsigned(1023, AMPLITUDE_WIDTH),
 998 => to_unsigned(1023, AMPLITUDE_WIDTH),
 999 => to_unsigned(1023, AMPLITUDE_WIDTH),
1000 => to_unsigned(1023, AMPLITUDE_WIDTH),
1001 => to_unsigned(1023, AMPLITUDE_WIDTH),
1002 => to_unsigned(1023, AMPLITUDE_WIDTH),
1003 => to_unsigned(1023, AMPLITUDE_WIDTH),
1004 => to_unsigned(1023, AMPLITUDE_WIDTH),
1005 => to_unsigned(1023, AMPLITUDE_WIDTH),
1006 => to_unsigned(1023, AMPLITUDE_WIDTH),
1007 => to_unsigned(1023, AMPLITUDE_WIDTH),
1008 => to_unsigned(1023, AMPLITUDE_WIDTH),
1009 => to_unsigned(1023, AMPLITUDE_WIDTH),
1010 => to_unsigned(1023, AMPLITUDE_WIDTH),
1011 => to_unsigned(1023, AMPLITUDE_WIDTH),
1012 => to_unsigned(1023, AMPLITUDE_WIDTH),
1013 => to_unsigned(1023, AMPLITUDE_WIDTH),
1014 => to_unsigned(1023, AMPLITUDE_WIDTH),
1015 => to_unsigned(1023, AMPLITUDE_WIDTH),
1016 => to_unsigned(1023, AMPLITUDE_WIDTH),
1017 => to_unsigned(1023, AMPLITUDE_WIDTH),
1018 => to_unsigned(1023, AMPLITUDE_WIDTH),
1019 => to_unsigned(1023, AMPLITUDE_WIDTH),
1020 => to_unsigned(1023, AMPLITUDE_WIDTH),
1021 => to_unsigned(1023, AMPLITUDE_WIDTH),
1022 => to_unsigned(1023, AMPLITUDE_WIDTH),
1023 => to_unsigned(1023, AMPLITUDE_WIDTH)
);
    
end lut_pkg;