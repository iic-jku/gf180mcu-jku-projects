module phase_to_amplitude
  (input  clock_i,
   input  reset_i,
   input  [31:0] phase_i,
   output [9:0] amplitude_o);
  wire [31:0] phase_reg;
  wire [31:0] phase_next;
  wire [11:0] address_reg;
  wire [11:0] address_next;
  wire [9:0] amplitude_reg;
  wire [9:0] amplitude_next;
  wire [11:0] n914;
  wire n916;
  wire n917;
  wire [9:0] n918;
  wire [9:0] n919;
  wire [9:0] n920;
  wire [9:0] n921;
  wire n928;
  wire n929;
  wire [9:0] n930;
  wire [9:0] n932;
  wire [9:0] n933;
  reg [31:0] n947;
  reg [11:0] n948;
  reg [9:0] n949;
  wire [9:0] n952; // mem_rd
  assign amplitude_o = amplitude_reg; //(module output)
  /* ../../vhdl/src/phase_to_amplitude.vhd:17:12  */
  assign phase_reg = n947; // (signal)
  /* ../../vhdl/src/phase_to_amplitude.vhd:18:12  */
  assign phase_next = phase_i; // (signal)
  /* ../../vhdl/src/phase_to_amplitude.vhd:19:12  */
  assign address_reg = n948; // (signal)
  /* ../../vhdl/src/phase_to_amplitude.vhd:20:12  */
  assign address_next = n914; // (signal)
  /* ../../vhdl/src/phase_to_amplitude.vhd:21:12  */
  assign amplitude_reg = n949; // (signal)
  /* ../../vhdl/src/phase_to_amplitude.vhd:22:12  */
  assign amplitude_next = n933; // (signal)
  /* ../../vhdl/src/phase_to_amplitude.vhd:37:34  */
  assign n914 = phase_reg[31:20]; // extract
  /* ../../vhdl/src/phase_to_amplitude.vhd:41:20  */
  assign n916 = address_reg[10]; // extract
  /* ../../vhdl/src/phase_to_amplitude.vhd:41:24  */
  assign n917 = ~n916;
  /* ../../vhdl/src/phase_to_amplitude.vhd:42:39  */
  assign n918 = address_reg[9:0]; // extract
  /* ../../vhdl/src/phase_to_amplitude.vhd:44:43  */
  assign n919 = address_reg[9:0]; // extract
  /* ../../vhdl/src/phase_to_amplitude.vhd:44:28  */
  assign n920 = ~n919;
  /* ../../vhdl/src/phase_to_amplitude.vhd:41:9  */
  assign n921 = n917 ? n918 : n920;
  /* ../../vhdl/src/phase_to_amplitude.vhd:49:21  */
  assign n928 = address_reg[11]; // extract
  /* ../../vhdl/src/phase_to_amplitude.vhd:49:25  */
  assign n929 = ~n928;
  /* ../../vhdl/src/phase_to_amplitude.vhd:52:32  */
  assign n930 = ~n952;
  /* ../../vhdl/src/phase_to_amplitude.vhd:52:45  */
  assign n932 = n930 + 10'b0000000001;
  /* ../../vhdl/src/phase_to_amplitude.vhd:49:10  */
  assign n933 = n929 ? n952 : n932;
  /* ../../vhdl/src/phase_to_amplitude.vhd:62:9  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n947 <= 32'b00000000000000000000000000000000;
    else
      n947 <= phase_next;
  /* ../../vhdl/src/phase_to_amplitude.vhd:62:9  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n948 <= 12'b000000000000;
    else
      n948 <= address_next;
  /* ../../vhdl/src/phase_to_amplitude.vhd:62:9  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n949 <= 10'b0000000000;
    else
      n949 <= amplitude_next;
  /* ../../vhdl/src/phase_to_amplitude.vhd:47:28  */
  reg [9:0] n950[1023:0] ; // memory
  initial begin
    n950[1023] = 10'b1111111111;
    n950[1022] = 10'b1111111111;
    n950[1021] = 10'b1111111111;
    n950[1020] = 10'b1111111111;
    n950[1019] = 10'b1111111111;
    n950[1018] = 10'b1111111111;
    n950[1017] = 10'b1111111111;
    n950[1016] = 10'b1111111111;
    n950[1015] = 10'b1111111111;
    n950[1014] = 10'b1111111111;
    n950[1013] = 10'b1111111111;
    n950[1012] = 10'b1111111111;
    n950[1011] = 10'b1111111111;
    n950[1010] = 10'b1111111111;
    n950[1009] = 10'b1111111111;
    n950[1008] = 10'b1111111111;
    n950[1007] = 10'b1111111111;
    n950[1006] = 10'b1111111111;
    n950[1005] = 10'b1111111111;
    n950[1004] = 10'b1111111111;
    n950[1003] = 10'b1111111111;
    n950[1002] = 10'b1111111111;
    n950[1001] = 10'b1111111111;
    n950[1000] = 10'b1111111111;
    n950[999] = 10'b1111111111;
    n950[998] = 10'b1111111111;
    n950[997] = 10'b1111111111;
    n950[996] = 10'b1111111111;
    n950[995] = 10'b1111111111;
    n950[994] = 10'b1111111110;
    n950[993] = 10'b1111111110;
    n950[992] = 10'b1111111110;
    n950[991] = 10'b1111111110;
    n950[990] = 10'b1111111110;
    n950[989] = 10'b1111111110;
    n950[988] = 10'b1111111110;
    n950[987] = 10'b1111111110;
    n950[986] = 10'b1111111110;
    n950[985] = 10'b1111111110;
    n950[984] = 10'b1111111110;
    n950[983] = 10'b1111111110;
    n950[982] = 10'b1111111110;
    n950[981] = 10'b1111111110;
    n950[980] = 10'b1111111110;
    n950[979] = 10'b1111111110;
    n950[978] = 10'b1111111110;
    n950[977] = 10'b1111111110;
    n950[976] = 10'b1111111110;
    n950[975] = 10'b1111111110;
    n950[974] = 10'b1111111110;
    n950[973] = 10'b1111111101;
    n950[972] = 10'b1111111101;
    n950[971] = 10'b1111111101;
    n950[970] = 10'b1111111101;
    n950[969] = 10'b1111111101;
    n950[968] = 10'b1111111101;
    n950[967] = 10'b1111111101;
    n950[966] = 10'b1111111101;
    n950[965] = 10'b1111111101;
    n950[964] = 10'b1111111101;
    n950[963] = 10'b1111111101;
    n950[962] = 10'b1111111101;
    n950[961] = 10'b1111111101;
    n950[960] = 10'b1111111101;
    n950[959] = 10'b1111111101;
    n950[958] = 10'b1111111100;
    n950[957] = 10'b1111111100;
    n950[956] = 10'b1111111100;
    n950[955] = 10'b1111111100;
    n950[954] = 10'b1111111100;
    n950[953] = 10'b1111111100;
    n950[952] = 10'b1111111100;
    n950[951] = 10'b1111111100;
    n950[950] = 10'b1111111100;
    n950[949] = 10'b1111111100;
    n950[948] = 10'b1111111100;
    n950[947] = 10'b1111111100;
    n950[946] = 10'b1111111011;
    n950[945] = 10'b1111111011;
    n950[944] = 10'b1111111011;
    n950[943] = 10'b1111111011;
    n950[942] = 10'b1111111011;
    n950[941] = 10'b1111111011;
    n950[940] = 10'b1111111011;
    n950[939] = 10'b1111111011;
    n950[938] = 10'b1111111011;
    n950[937] = 10'b1111111011;
    n950[936] = 10'b1111111010;
    n950[935] = 10'b1111111010;
    n950[934] = 10'b1111111010;
    n950[933] = 10'b1111111010;
    n950[932] = 10'b1111111010;
    n950[931] = 10'b1111111010;
    n950[930] = 10'b1111111010;
    n950[929] = 10'b1111111010;
    n950[928] = 10'b1111111010;
    n950[927] = 10'b1111111001;
    n950[926] = 10'b1111111001;
    n950[925] = 10'b1111111001;
    n950[924] = 10'b1111111001;
    n950[923] = 10'b1111111001;
    n950[922] = 10'b1111111001;
    n950[921] = 10'b1111111001;
    n950[920] = 10'b1111111001;
    n950[919] = 10'b1111111000;
    n950[918] = 10'b1111111000;
    n950[917] = 10'b1111111000;
    n950[916] = 10'b1111111000;
    n950[915] = 10'b1111111000;
    n950[914] = 10'b1111111000;
    n950[913] = 10'b1111111000;
    n950[912] = 10'b1111111000;
    n950[911] = 10'b1111110111;
    n950[910] = 10'b1111110111;
    n950[909] = 10'b1111110111;
    n950[908] = 10'b1111110111;
    n950[907] = 10'b1111110111;
    n950[906] = 10'b1111110111;
    n950[905] = 10'b1111110111;
    n950[904] = 10'b1111110110;
    n950[903] = 10'b1111110110;
    n950[902] = 10'b1111110110;
    n950[901] = 10'b1111110110;
    n950[900] = 10'b1111110110;
    n950[899] = 10'b1111110110;
    n950[898] = 10'b1111110110;
    n950[897] = 10'b1111110101;
    n950[896] = 10'b1111110101;
    n950[895] = 10'b1111110101;
    n950[894] = 10'b1111110101;
    n950[893] = 10'b1111110101;
    n950[892] = 10'b1111110101;
    n950[891] = 10'b1111110101;
    n950[890] = 10'b1111110100;
    n950[889] = 10'b1111110100;
    n950[888] = 10'b1111110100;
    n950[887] = 10'b1111110100;
    n950[886] = 10'b1111110100;
    n950[885] = 10'b1111110100;
    n950[884] = 10'b1111110011;
    n950[883] = 10'b1111110011;
    n950[882] = 10'b1111110011;
    n950[881] = 10'b1111110011;
    n950[880] = 10'b1111110011;
    n950[879] = 10'b1111110011;
    n950[878] = 10'b1111110010;
    n950[877] = 10'b1111110010;
    n950[876] = 10'b1111110010;
    n950[875] = 10'b1111110010;
    n950[874] = 10'b1111110010;
    n950[873] = 10'b1111110001;
    n950[872] = 10'b1111110001;
    n950[871] = 10'b1111110001;
    n950[870] = 10'b1111110001;
    n950[869] = 10'b1111110001;
    n950[868] = 10'b1111110001;
    n950[867] = 10'b1111110000;
    n950[866] = 10'b1111110000;
    n950[865] = 10'b1111110000;
    n950[864] = 10'b1111110000;
    n950[863] = 10'b1111110000;
    n950[862] = 10'b1111101111;
    n950[861] = 10'b1111101111;
    n950[860] = 10'b1111101111;
    n950[859] = 10'b1111101111;
    n950[858] = 10'b1111101111;
    n950[857] = 10'b1111101110;
    n950[856] = 10'b1111101110;
    n950[855] = 10'b1111101110;
    n950[854] = 10'b1111101110;
    n950[853] = 10'b1111101110;
    n950[852] = 10'b1111101101;
    n950[851] = 10'b1111101101;
    n950[850] = 10'b1111101101;
    n950[849] = 10'b1111101101;
    n950[848] = 10'b1111101101;
    n950[847] = 10'b1111101100;
    n950[846] = 10'b1111101100;
    n950[845] = 10'b1111101100;
    n950[844] = 10'b1111101100;
    n950[843] = 10'b1111101100;
    n950[842] = 10'b1111101011;
    n950[841] = 10'b1111101011;
    n950[840] = 10'b1111101011;
    n950[839] = 10'b1111101011;
    n950[838] = 10'b1111101011;
    n950[837] = 10'b1111101010;
    n950[836] = 10'b1111101010;
    n950[835] = 10'b1111101010;
    n950[834] = 10'b1111101010;
    n950[833] = 10'b1111101001;
    n950[832] = 10'b1111101001;
    n950[831] = 10'b1111101001;
    n950[830] = 10'b1111101001;
    n950[829] = 10'b1111101000;
    n950[828] = 10'b1111101000;
    n950[827] = 10'b1111101000;
    n950[826] = 10'b1111101000;
    n950[825] = 10'b1111101000;
    n950[824] = 10'b1111100111;
    n950[823] = 10'b1111100111;
    n950[822] = 10'b1111100111;
    n950[821] = 10'b1111100111;
    n950[820] = 10'b1111100110;
    n950[819] = 10'b1111100110;
    n950[818] = 10'b1111100110;
    n950[817] = 10'b1111100110;
    n950[816] = 10'b1111100101;
    n950[815] = 10'b1111100101;
    n950[814] = 10'b1111100101;
    n950[813] = 10'b1111100101;
    n950[812] = 10'b1111100100;
    n950[811] = 10'b1111100100;
    n950[810] = 10'b1111100100;
    n950[809] = 10'b1111100100;
    n950[808] = 10'b1111100011;
    n950[807] = 10'b1111100011;
    n950[806] = 10'b1111100011;
    n950[805] = 10'b1111100011;
    n950[804] = 10'b1111100010;
    n950[803] = 10'b1111100010;
    n950[802] = 10'b1111100010;
    n950[801] = 10'b1111100010;
    n950[800] = 10'b1111100001;
    n950[799] = 10'b1111100001;
    n950[798] = 10'b1111100001;
    n950[797] = 10'b1111100001;
    n950[796] = 10'b1111100000;
    n950[795] = 10'b1111100000;
    n950[794] = 10'b1111100000;
    n950[793] = 10'b1111011111;
    n950[792] = 10'b1111011111;
    n950[791] = 10'b1111011111;
    n950[790] = 10'b1111011111;
    n950[789] = 10'b1111011110;
    n950[788] = 10'b1111011110;
    n950[787] = 10'b1111011110;
    n950[786] = 10'b1111011110;
    n950[785] = 10'b1111011101;
    n950[784] = 10'b1111011101;
    n950[783] = 10'b1111011101;
    n950[782] = 10'b1111011100;
    n950[781] = 10'b1111011100;
    n950[780] = 10'b1111011100;
    n950[779] = 10'b1111011100;
    n950[778] = 10'b1111011011;
    n950[777] = 10'b1111011011;
    n950[776] = 10'b1111011011;
    n950[775] = 10'b1111011010;
    n950[774] = 10'b1111011010;
    n950[773] = 10'b1111011010;
    n950[772] = 10'b1111011001;
    n950[771] = 10'b1111011001;
    n950[770] = 10'b1111011001;
    n950[769] = 10'b1111011001;
    n950[768] = 10'b1111011000;
    n950[767] = 10'b1111011000;
    n950[766] = 10'b1111011000;
    n950[765] = 10'b1111010111;
    n950[764] = 10'b1111010111;
    n950[763] = 10'b1111010111;
    n950[762] = 10'b1111010110;
    n950[761] = 10'b1111010110;
    n950[760] = 10'b1111010110;
    n950[759] = 10'b1111010110;
    n950[758] = 10'b1111010101;
    n950[757] = 10'b1111010101;
    n950[756] = 10'b1111010101;
    n950[755] = 10'b1111010100;
    n950[754] = 10'b1111010100;
    n950[753] = 10'b1111010100;
    n950[752] = 10'b1111010011;
    n950[751] = 10'b1111010011;
    n950[750] = 10'b1111010011;
    n950[749] = 10'b1111010010;
    n950[748] = 10'b1111010010;
    n950[747] = 10'b1111010010;
    n950[746] = 10'b1111010001;
    n950[745] = 10'b1111010001;
    n950[744] = 10'b1111010001;
    n950[743] = 10'b1111010000;
    n950[742] = 10'b1111010000;
    n950[741] = 10'b1111010000;
    n950[740] = 10'b1111001111;
    n950[739] = 10'b1111001111;
    n950[738] = 10'b1111001111;
    n950[737] = 10'b1111001110;
    n950[736] = 10'b1111001110;
    n950[735] = 10'b1111001110;
    n950[734] = 10'b1111001101;
    n950[733] = 10'b1111001101;
    n950[732] = 10'b1111001101;
    n950[731] = 10'b1111001100;
    n950[730] = 10'b1111001100;
    n950[729] = 10'b1111001100;
    n950[728] = 10'b1111001011;
    n950[727] = 10'b1111001011;
    n950[726] = 10'b1111001011;
    n950[725] = 10'b1111001010;
    n950[724] = 10'b1111001010;
    n950[723] = 10'b1111001010;
    n950[722] = 10'b1111001001;
    n950[721] = 10'b1111001001;
    n950[720] = 10'b1111001001;
    n950[719] = 10'b1111001000;
    n950[718] = 10'b1111001000;
    n950[717] = 10'b1111001000;
    n950[716] = 10'b1111000111;
    n950[715] = 10'b1111000111;
    n950[714] = 10'b1111000110;
    n950[713] = 10'b1111000110;
    n950[712] = 10'b1111000110;
    n950[711] = 10'b1111000101;
    n950[710] = 10'b1111000101;
    n950[709] = 10'b1111000101;
    n950[708] = 10'b1111000100;
    n950[707] = 10'b1111000100;
    n950[706] = 10'b1111000100;
    n950[705] = 10'b1111000011;
    n950[704] = 10'b1111000011;
    n950[703] = 10'b1111000010;
    n950[702] = 10'b1111000010;
    n950[701] = 10'b1111000010;
    n950[700] = 10'b1111000001;
    n950[699] = 10'b1111000001;
    n950[698] = 10'b1111000001;
    n950[697] = 10'b1111000000;
    n950[696] = 10'b1111000000;
    n950[695] = 10'b1110111111;
    n950[694] = 10'b1110111111;
    n950[693] = 10'b1110111111;
    n950[692] = 10'b1110111110;
    n950[691] = 10'b1110111110;
    n950[690] = 10'b1110111110;
    n950[689] = 10'b1110111101;
    n950[688] = 10'b1110111101;
    n950[687] = 10'b1110111100;
    n950[686] = 10'b1110111100;
    n950[685] = 10'b1110111100;
    n950[684] = 10'b1110111011;
    n950[683] = 10'b1110111011;
    n950[682] = 10'b1110111010;
    n950[681] = 10'b1110111010;
    n950[680] = 10'b1110111010;
    n950[679] = 10'b1110111001;
    n950[678] = 10'b1110111001;
    n950[677] = 10'b1110111000;
    n950[676] = 10'b1110111000;
    n950[675] = 10'b1110111000;
    n950[674] = 10'b1110110111;
    n950[673] = 10'b1110110111;
    n950[672] = 10'b1110110110;
    n950[671] = 10'b1110110110;
    n950[670] = 10'b1110110110;
    n950[669] = 10'b1110110101;
    n950[668] = 10'b1110110101;
    n950[667] = 10'b1110110100;
    n950[666] = 10'b1110110100;
    n950[665] = 10'b1110110100;
    n950[664] = 10'b1110110011;
    n950[663] = 10'b1110110011;
    n950[662] = 10'b1110110010;
    n950[661] = 10'b1110110010;
    n950[660] = 10'b1110110010;
    n950[659] = 10'b1110110001;
    n950[658] = 10'b1110110001;
    n950[657] = 10'b1110110000;
    n950[656] = 10'b1110110000;
    n950[655] = 10'b1110101111;
    n950[654] = 10'b1110101111;
    n950[653] = 10'b1110101111;
    n950[652] = 10'b1110101110;
    n950[651] = 10'b1110101110;
    n950[650] = 10'b1110101101;
    n950[649] = 10'b1110101101;
    n950[648] = 10'b1110101101;
    n950[647] = 10'b1110101100;
    n950[646] = 10'b1110101100;
    n950[645] = 10'b1110101011;
    n950[644] = 10'b1110101011;
    n950[643] = 10'b1110101010;
    n950[642] = 10'b1110101010;
    n950[641] = 10'b1110101010;
    n950[640] = 10'b1110101001;
    n950[639] = 10'b1110101001;
    n950[638] = 10'b1110101000;
    n950[637] = 10'b1110101000;
    n950[636] = 10'b1110100111;
    n950[635] = 10'b1110100111;
    n950[634] = 10'b1110100110;
    n950[633] = 10'b1110100110;
    n950[632] = 10'b1110100110;
    n950[631] = 10'b1110100101;
    n950[630] = 10'b1110100101;
    n950[629] = 10'b1110100100;
    n950[628] = 10'b1110100100;
    n950[627] = 10'b1110100011;
    n950[626] = 10'b1110100011;
    n950[625] = 10'b1110100010;
    n950[624] = 10'b1110100010;
    n950[623] = 10'b1110100010;
    n950[622] = 10'b1110100001;
    n950[621] = 10'b1110100001;
    n950[620] = 10'b1110100000;
    n950[619] = 10'b1110100000;
    n950[618] = 10'b1110011111;
    n950[617] = 10'b1110011111;
    n950[616] = 10'b1110011110;
    n950[615] = 10'b1110011110;
    n950[614] = 10'b1110011101;
    n950[613] = 10'b1110011101;
    n950[612] = 10'b1110011100;
    n950[611] = 10'b1110011100;
    n950[610] = 10'b1110011100;
    n950[609] = 10'b1110011011;
    n950[608] = 10'b1110011011;
    n950[607] = 10'b1110011010;
    n950[606] = 10'b1110011010;
    n950[605] = 10'b1110011001;
    n950[604] = 10'b1110011001;
    n950[603] = 10'b1110011000;
    n950[602] = 10'b1110011000;
    n950[601] = 10'b1110010111;
    n950[600] = 10'b1110010111;
    n950[599] = 10'b1110010110;
    n950[598] = 10'b1110010110;
    n950[597] = 10'b1110010101;
    n950[596] = 10'b1110010101;
    n950[595] = 10'b1110010100;
    n950[594] = 10'b1110010100;
    n950[593] = 10'b1110010100;
    n950[592] = 10'b1110010011;
    n950[591] = 10'b1110010011;
    n950[590] = 10'b1110010010;
    n950[589] = 10'b1110010010;
    n950[588] = 10'b1110010001;
    n950[587] = 10'b1110010001;
    n950[586] = 10'b1110010000;
    n950[585] = 10'b1110010000;
    n950[584] = 10'b1110001111;
    n950[583] = 10'b1110001111;
    n950[582] = 10'b1110001110;
    n950[581] = 10'b1110001110;
    n950[580] = 10'b1110001101;
    n950[579] = 10'b1110001101;
    n950[578] = 10'b1110001100;
    n950[577] = 10'b1110001100;
    n950[576] = 10'b1110001011;
    n950[575] = 10'b1110001011;
    n950[574] = 10'b1110001010;
    n950[573] = 10'b1110001010;
    n950[572] = 10'b1110001001;
    n950[571] = 10'b1110001001;
    n950[570] = 10'b1110001000;
    n950[569] = 10'b1110001000;
    n950[568] = 10'b1110000111;
    n950[567] = 10'b1110000111;
    n950[566] = 10'b1110000110;
    n950[565] = 10'b1110000110;
    n950[564] = 10'b1110000101;
    n950[563] = 10'b1110000101;
    n950[562] = 10'b1110000100;
    n950[561] = 10'b1110000100;
    n950[560] = 10'b1110000011;
    n950[559] = 10'b1110000011;
    n950[558] = 10'b1110000010;
    n950[557] = 10'b1110000010;
    n950[556] = 10'b1110000001;
    n950[555] = 10'b1110000001;
    n950[554] = 10'b1110000000;
    n950[553] = 10'b1101111111;
    n950[552] = 10'b1101111111;
    n950[551] = 10'b1101111110;
    n950[550] = 10'b1101111110;
    n950[549] = 10'b1101111101;
    n950[548] = 10'b1101111101;
    n950[547] = 10'b1101111100;
    n950[546] = 10'b1101111100;
    n950[545] = 10'b1101111011;
    n950[544] = 10'b1101111011;
    n950[543] = 10'b1101111010;
    n950[542] = 10'b1101111010;
    n950[541] = 10'b1101111001;
    n950[540] = 10'b1101111001;
    n950[539] = 10'b1101111000;
    n950[538] = 10'b1101111000;
    n950[537] = 10'b1101110111;
    n950[536] = 10'b1101110111;
    n950[535] = 10'b1101110110;
    n950[534] = 10'b1101110101;
    n950[533] = 10'b1101110101;
    n950[532] = 10'b1101110100;
    n950[531] = 10'b1101110100;
    n950[530] = 10'b1101110011;
    n950[529] = 10'b1101110011;
    n950[528] = 10'b1101110010;
    n950[527] = 10'b1101110010;
    n950[526] = 10'b1101110001;
    n950[525] = 10'b1101110001;
    n950[524] = 10'b1101110000;
    n950[523] = 10'b1101110000;
    n950[522] = 10'b1101101111;
    n950[521] = 10'b1101101110;
    n950[520] = 10'b1101101110;
    n950[519] = 10'b1101101101;
    n950[518] = 10'b1101101101;
    n950[517] = 10'b1101101100;
    n950[516] = 10'b1101101100;
    n950[515] = 10'b1101101011;
    n950[514] = 10'b1101101011;
    n950[513] = 10'b1101101010;
    n950[512] = 10'b1101101001;
    n950[511] = 10'b1101101001;
    n950[510] = 10'b1101101000;
    n950[509] = 10'b1101101000;
    n950[508] = 10'b1101100111;
    n950[507] = 10'b1101100111;
    n950[506] = 10'b1101100110;
    n950[505] = 10'b1101100110;
    n950[504] = 10'b1101100101;
    n950[503] = 10'b1101100100;
    n950[502] = 10'b1101100100;
    n950[501] = 10'b1101100011;
    n950[500] = 10'b1101100011;
    n950[499] = 10'b1101100010;
    n950[498] = 10'b1101100010;
    n950[497] = 10'b1101100001;
    n950[496] = 10'b1101100000;
    n950[495] = 10'b1101100000;
    n950[494] = 10'b1101011111;
    n950[493] = 10'b1101011111;
    n950[492] = 10'b1101011110;
    n950[491] = 10'b1101011110;
    n950[490] = 10'b1101011101;
    n950[489] = 10'b1101011100;
    n950[488] = 10'b1101011100;
    n950[487] = 10'b1101011011;
    n950[486] = 10'b1101011011;
    n950[485] = 10'b1101011010;
    n950[484] = 10'b1101011010;
    n950[483] = 10'b1101011001;
    n950[482] = 10'b1101011000;
    n950[481] = 10'b1101011000;
    n950[480] = 10'b1101010111;
    n950[479] = 10'b1101010111;
    n950[478] = 10'b1101010110;
    n950[477] = 10'b1101010110;
    n950[476] = 10'b1101010101;
    n950[475] = 10'b1101010100;
    n950[474] = 10'b1101010100;
    n950[473] = 10'b1101010011;
    n950[472] = 10'b1101010011;
    n950[471] = 10'b1101010010;
    n950[470] = 10'b1101010001;
    n950[469] = 10'b1101010001;
    n950[468] = 10'b1101010000;
    n950[467] = 10'b1101010000;
    n950[466] = 10'b1101001111;
    n950[465] = 10'b1101001110;
    n950[464] = 10'b1101001110;
    n950[463] = 10'b1101001101;
    n950[462] = 10'b1101001101;
    n950[461] = 10'b1101001100;
    n950[460] = 10'b1101001011;
    n950[459] = 10'b1101001011;
    n950[458] = 10'b1101001010;
    n950[457] = 10'b1101001010;
    n950[456] = 10'b1101001001;
    n950[455] = 10'b1101001000;
    n950[454] = 10'b1101001000;
    n950[453] = 10'b1101000111;
    n950[452] = 10'b1101000111;
    n950[451] = 10'b1101000110;
    n950[450] = 10'b1101000101;
    n950[449] = 10'b1101000101;
    n950[448] = 10'b1101000100;
    n950[447] = 10'b1101000100;
    n950[446] = 10'b1101000011;
    n950[445] = 10'b1101000010;
    n950[444] = 10'b1101000010;
    n950[443] = 10'b1101000001;
    n950[442] = 10'b1101000001;
    n950[441] = 10'b1101000000;
    n950[440] = 10'b1100111111;
    n950[439] = 10'b1100111111;
    n950[438] = 10'b1100111110;
    n950[437] = 10'b1100111110;
    n950[436] = 10'b1100111101;
    n950[435] = 10'b1100111100;
    n950[434] = 10'b1100111100;
    n950[433] = 10'b1100111011;
    n950[432] = 10'b1100111010;
    n950[431] = 10'b1100111010;
    n950[430] = 10'b1100111001;
    n950[429] = 10'b1100111001;
    n950[428] = 10'b1100111000;
    n950[427] = 10'b1100110111;
    n950[426] = 10'b1100110111;
    n950[425] = 10'b1100110110;
    n950[424] = 10'b1100110101;
    n950[423] = 10'b1100110101;
    n950[422] = 10'b1100110100;
    n950[421] = 10'b1100110100;
    n950[420] = 10'b1100110011;
    n950[419] = 10'b1100110010;
    n950[418] = 10'b1100110010;
    n950[417] = 10'b1100110001;
    n950[416] = 10'b1100110000;
    n950[415] = 10'b1100110000;
    n950[414] = 10'b1100101111;
    n950[413] = 10'b1100101111;
    n950[412] = 10'b1100101110;
    n950[411] = 10'b1100101101;
    n950[410] = 10'b1100101101;
    n950[409] = 10'b1100101100;
    n950[408] = 10'b1100101011;
    n950[407] = 10'b1100101011;
    n950[406] = 10'b1100101010;
    n950[405] = 10'b1100101001;
    n950[404] = 10'b1100101001;
    n950[403] = 10'b1100101000;
    n950[402] = 10'b1100101000;
    n950[401] = 10'b1100100111;
    n950[400] = 10'b1100100110;
    n950[399] = 10'b1100100110;
    n950[398] = 10'b1100100101;
    n950[397] = 10'b1100100100;
    n950[396] = 10'b1100100100;
    n950[395] = 10'b1100100011;
    n950[394] = 10'b1100100010;
    n950[393] = 10'b1100100010;
    n950[392] = 10'b1100100001;
    n950[391] = 10'b1100100000;
    n950[390] = 10'b1100100000;
    n950[389] = 10'b1100011111;
    n950[388] = 10'b1100011111;
    n950[387] = 10'b1100011110;
    n950[386] = 10'b1100011101;
    n950[385] = 10'b1100011101;
    n950[384] = 10'b1100011100;
    n950[383] = 10'b1100011011;
    n950[382] = 10'b1100011011;
    n950[381] = 10'b1100011010;
    n950[380] = 10'b1100011001;
    n950[379] = 10'b1100011001;
    n950[378] = 10'b1100011000;
    n950[377] = 10'b1100010111;
    n950[376] = 10'b1100010111;
    n950[375] = 10'b1100010110;
    n950[374] = 10'b1100010101;
    n950[373] = 10'b1100010101;
    n950[372] = 10'b1100010100;
    n950[371] = 10'b1100010011;
    n950[370] = 10'b1100010011;
    n950[369] = 10'b1100010010;
    n950[368] = 10'b1100010001;
    n950[367] = 10'b1100010001;
    n950[366] = 10'b1100010000;
    n950[365] = 10'b1100001111;
    n950[364] = 10'b1100001111;
    n950[363] = 10'b1100001110;
    n950[362] = 10'b1100001101;
    n950[361] = 10'b1100001101;
    n950[360] = 10'b1100001100;
    n950[359] = 10'b1100001011;
    n950[358] = 10'b1100001011;
    n950[357] = 10'b1100001010;
    n950[356] = 10'b1100001001;
    n950[355] = 10'b1100001001;
    n950[354] = 10'b1100001000;
    n950[353] = 10'b1100000111;
    n950[352] = 10'b1100000111;
    n950[351] = 10'b1100000110;
    n950[350] = 10'b1100000101;
    n950[349] = 10'b1100000101;
    n950[348] = 10'b1100000100;
    n950[347] = 10'b1100000011;
    n950[346] = 10'b1100000011;
    n950[345] = 10'b1100000010;
    n950[344] = 10'b1100000001;
    n950[343] = 10'b1100000001;
    n950[342] = 10'b1100000000;
    n950[341] = 10'b1011111111;
    n950[340] = 10'b1011111111;
    n950[339] = 10'b1011111110;
    n950[338] = 10'b1011111101;
    n950[337] = 10'b1011111101;
    n950[336] = 10'b1011111100;
    n950[335] = 10'b1011111011;
    n950[334] = 10'b1011111010;
    n950[333] = 10'b1011111010;
    n950[332] = 10'b1011111001;
    n950[331] = 10'b1011111000;
    n950[330] = 10'b1011111000;
    n950[329] = 10'b1011110111;
    n950[328] = 10'b1011110110;
    n950[327] = 10'b1011110110;
    n950[326] = 10'b1011110101;
    n950[325] = 10'b1011110100;
    n950[324] = 10'b1011110100;
    n950[323] = 10'b1011110011;
    n950[322] = 10'b1011110010;
    n950[321] = 10'b1011110010;
    n950[320] = 10'b1011110001;
    n950[319] = 10'b1011110000;
    n950[318] = 10'b1011101111;
    n950[317] = 10'b1011101111;
    n950[316] = 10'b1011101110;
    n950[315] = 10'b1011101101;
    n950[314] = 10'b1011101101;
    n950[313] = 10'b1011101100;
    n950[312] = 10'b1011101011;
    n950[311] = 10'b1011101011;
    n950[310] = 10'b1011101010;
    n950[309] = 10'b1011101001;
    n950[308] = 10'b1011101000;
    n950[307] = 10'b1011101000;
    n950[306] = 10'b1011100111;
    n950[305] = 10'b1011100110;
    n950[304] = 10'b1011100110;
    n950[303] = 10'b1011100101;
    n950[302] = 10'b1011100100;
    n950[301] = 10'b1011100100;
    n950[300] = 10'b1011100011;
    n950[299] = 10'b1011100010;
    n950[298] = 10'b1011100001;
    n950[297] = 10'b1011100001;
    n950[296] = 10'b1011100000;
    n950[295] = 10'b1011011111;
    n950[294] = 10'b1011011111;
    n950[293] = 10'b1011011110;
    n950[292] = 10'b1011011101;
    n950[291] = 10'b1011011101;
    n950[290] = 10'b1011011100;
    n950[289] = 10'b1011011011;
    n950[288] = 10'b1011011010;
    n950[287] = 10'b1011011010;
    n950[286] = 10'b1011011001;
    n950[285] = 10'b1011011000;
    n950[284] = 10'b1011011000;
    n950[283] = 10'b1011010111;
    n950[282] = 10'b1011010110;
    n950[281] = 10'b1011010101;
    n950[280] = 10'b1011010101;
    n950[279] = 10'b1011010100;
    n950[278] = 10'b1011010011;
    n950[277] = 10'b1011010011;
    n950[276] = 10'b1011010010;
    n950[275] = 10'b1011010001;
    n950[274] = 10'b1011010000;
    n950[273] = 10'b1011010000;
    n950[272] = 10'b1011001111;
    n950[271] = 10'b1011001110;
    n950[270] = 10'b1011001110;
    n950[269] = 10'b1011001101;
    n950[268] = 10'b1011001100;
    n950[267] = 10'b1011001011;
    n950[266] = 10'b1011001011;
    n950[265] = 10'b1011001010;
    n950[264] = 10'b1011001001;
    n950[263] = 10'b1011001000;
    n950[262] = 10'b1011001000;
    n950[261] = 10'b1011000111;
    n950[260] = 10'b1011000110;
    n950[259] = 10'b1011000110;
    n950[258] = 10'b1011000101;
    n950[257] = 10'b1011000100;
    n950[256] = 10'b1011000011;
    n950[255] = 10'b1011000011;
    n950[254] = 10'b1011000010;
    n950[253] = 10'b1011000001;
    n950[252] = 10'b1011000001;
    n950[251] = 10'b1011000000;
    n950[250] = 10'b1010111111;
    n950[249] = 10'b1010111110;
    n950[248] = 10'b1010111110;
    n950[247] = 10'b1010111101;
    n950[246] = 10'b1010111100;
    n950[245] = 10'b1010111011;
    n950[244] = 10'b1010111011;
    n950[243] = 10'b1010111010;
    n950[242] = 10'b1010111001;
    n950[241] = 10'b1010111000;
    n950[240] = 10'b1010111000;
    n950[239] = 10'b1010110111;
    n950[238] = 10'b1010110110;
    n950[237] = 10'b1010110110;
    n950[236] = 10'b1010110101;
    n950[235] = 10'b1010110100;
    n950[234] = 10'b1010110011;
    n950[233] = 10'b1010110011;
    n950[232] = 10'b1010110010;
    n950[231] = 10'b1010110001;
    n950[230] = 10'b1010110000;
    n950[229] = 10'b1010110000;
    n950[228] = 10'b1010101111;
    n950[227] = 10'b1010101110;
    n950[226] = 10'b1010101101;
    n950[225] = 10'b1010101101;
    n950[224] = 10'b1010101100;
    n950[223] = 10'b1010101011;
    n950[222] = 10'b1010101011;
    n950[221] = 10'b1010101010;
    n950[220] = 10'b1010101001;
    n950[219] = 10'b1010101000;
    n950[218] = 10'b1010101000;
    n950[217] = 10'b1010100111;
    n950[216] = 10'b1010100110;
    n950[215] = 10'b1010100101;
    n950[214] = 10'b1010100101;
    n950[213] = 10'b1010100100;
    n950[212] = 10'b1010100011;
    n950[211] = 10'b1010100010;
    n950[210] = 10'b1010100010;
    n950[209] = 10'b1010100001;
    n950[208] = 10'b1010100000;
    n950[207] = 10'b1010011111;
    n950[206] = 10'b1010011111;
    n950[205] = 10'b1010011110;
    n950[204] = 10'b1010011101;
    n950[203] = 10'b1010011100;
    n950[202] = 10'b1010011100;
    n950[201] = 10'b1010011011;
    n950[200] = 10'b1010011010;
    n950[199] = 10'b1010011001;
    n950[198] = 10'b1010011001;
    n950[197] = 10'b1010011000;
    n950[196] = 10'b1010010111;
    n950[195] = 10'b1010010110;
    n950[194] = 10'b1010010110;
    n950[193] = 10'b1010010101;
    n950[192] = 10'b1010010100;
    n950[191] = 10'b1010010011;
    n950[190] = 10'b1010010011;
    n950[189] = 10'b1010010010;
    n950[188] = 10'b1010010001;
    n950[187] = 10'b1010010000;
    n950[186] = 10'b1010010000;
    n950[185] = 10'b1010001111;
    n950[184] = 10'b1010001110;
    n950[183] = 10'b1010001101;
    n950[182] = 10'b1010001101;
    n950[181] = 10'b1010001100;
    n950[180] = 10'b1010001011;
    n950[179] = 10'b1010001010;
    n950[178] = 10'b1010001010;
    n950[177] = 10'b1010001001;
    n950[176] = 10'b1010001000;
    n950[175] = 10'b1010000111;
    n950[174] = 10'b1010000111;
    n950[173] = 10'b1010000110;
    n950[172] = 10'b1010000101;
    n950[171] = 10'b1010000100;
    n950[170] = 10'b1010000100;
    n950[169] = 10'b1010000011;
    n950[168] = 10'b1010000010;
    n950[167] = 10'b1010000001;
    n950[166] = 10'b1010000000;
    n950[165] = 10'b1010000000;
    n950[164] = 10'b1001111111;
    n950[163] = 10'b1001111110;
    n950[162] = 10'b1001111101;
    n950[161] = 10'b1001111101;
    n950[160] = 10'b1001111100;
    n950[159] = 10'b1001111011;
    n950[158] = 10'b1001111010;
    n950[157] = 10'b1001111010;
    n950[156] = 10'b1001111001;
    n950[155] = 10'b1001111000;
    n950[154] = 10'b1001110111;
    n950[153] = 10'b1001110111;
    n950[152] = 10'b1001110110;
    n950[151] = 10'b1001110101;
    n950[150] = 10'b1001110100;
    n950[149] = 10'b1001110100;
    n950[148] = 10'b1001110011;
    n950[147] = 10'b1001110010;
    n950[146] = 10'b1001110001;
    n950[145] = 10'b1001110000;
    n950[144] = 10'b1001110000;
    n950[143] = 10'b1001101111;
    n950[142] = 10'b1001101110;
    n950[141] = 10'b1001101101;
    n950[140] = 10'b1001101101;
    n950[139] = 10'b1001101100;
    n950[138] = 10'b1001101011;
    n950[137] = 10'b1001101010;
    n950[136] = 10'b1001101010;
    n950[135] = 10'b1001101001;
    n950[134] = 10'b1001101000;
    n950[133] = 10'b1001100111;
    n950[132] = 10'b1001100110;
    n950[131] = 10'b1001100110;
    n950[130] = 10'b1001100101;
    n950[129] = 10'b1001100100;
    n950[128] = 10'b1001100011;
    n950[127] = 10'b1001100011;
    n950[126] = 10'b1001100010;
    n950[125] = 10'b1001100001;
    n950[124] = 10'b1001100000;
    n950[123] = 10'b1001100000;
    n950[122] = 10'b1001011111;
    n950[121] = 10'b1001011110;
    n950[120] = 10'b1001011101;
    n950[119] = 10'b1001011100;
    n950[118] = 10'b1001011100;
    n950[117] = 10'b1001011011;
    n950[116] = 10'b1001011010;
    n950[115] = 10'b1001011001;
    n950[114] = 10'b1001011001;
    n950[113] = 10'b1001011000;
    n950[112] = 10'b1001010111;
    n950[111] = 10'b1001010110;
    n950[110] = 10'b1001010101;
    n950[109] = 10'b1001010101;
    n950[108] = 10'b1001010100;
    n950[107] = 10'b1001010011;
    n950[106] = 10'b1001010010;
    n950[105] = 10'b1001010010;
    n950[104] = 10'b1001010001;
    n950[103] = 10'b1001010000;
    n950[102] = 10'b1001001111;
    n950[101] = 10'b1001001111;
    n950[100] = 10'b1001001110;
    n950[99] = 10'b1001001101;
    n950[98] = 10'b1001001100;
    n950[97] = 10'b1001001011;
    n950[96] = 10'b1001001011;
    n950[95] = 10'b1001001010;
    n950[94] = 10'b1001001001;
    n950[93] = 10'b1001001000;
    n950[92] = 10'b1001001000;
    n950[91] = 10'b1001000111;
    n950[90] = 10'b1001000110;
    n950[89] = 10'b1001000101;
    n950[88] = 10'b1001000100;
    n950[87] = 10'b1001000100;
    n950[86] = 10'b1001000011;
    n950[85] = 10'b1001000010;
    n950[84] = 10'b1001000001;
    n950[83] = 10'b1001000001;
    n950[82] = 10'b1001000000;
    n950[81] = 10'b1000111111;
    n950[80] = 10'b1000111110;
    n950[79] = 10'b1000111101;
    n950[78] = 10'b1000111101;
    n950[77] = 10'b1000111100;
    n950[76] = 10'b1000111011;
    n950[75] = 10'b1000111010;
    n950[74] = 10'b1000111001;
    n950[73] = 10'b1000111001;
    n950[72] = 10'b1000111000;
    n950[71] = 10'b1000110111;
    n950[70] = 10'b1000110110;
    n950[69] = 10'b1000110110;
    n950[68] = 10'b1000110101;
    n950[67] = 10'b1000110100;
    n950[66] = 10'b1000110011;
    n950[65] = 10'b1000110010;
    n950[64] = 10'b1000110010;
    n950[63] = 10'b1000110001;
    n950[62] = 10'b1000110000;
    n950[61] = 10'b1000101111;
    n950[60] = 10'b1000101111;
    n950[59] = 10'b1000101110;
    n950[58] = 10'b1000101101;
    n950[57] = 10'b1000101100;
    n950[56] = 10'b1000101011;
    n950[55] = 10'b1000101011;
    n950[54] = 10'b1000101010;
    n950[53] = 10'b1000101001;
    n950[52] = 10'b1000101000;
    n950[51] = 10'b1000101000;
    n950[50] = 10'b1000100111;
    n950[49] = 10'b1000100110;
    n950[48] = 10'b1000100101;
    n950[47] = 10'b1000100100;
    n950[46] = 10'b1000100100;
    n950[45] = 10'b1000100011;
    n950[44] = 10'b1000100010;
    n950[43] = 10'b1000100001;
    n950[42] = 10'b1000100000;
    n950[41] = 10'b1000100000;
    n950[40] = 10'b1000011111;
    n950[39] = 10'b1000011110;
    n950[38] = 10'b1000011101;
    n950[37] = 10'b1000011101;
    n950[36] = 10'b1000011100;
    n950[35] = 10'b1000011011;
    n950[34] = 10'b1000011010;
    n950[33] = 10'b1000011001;
    n950[32] = 10'b1000011001;
    n950[31] = 10'b1000011000;
    n950[30] = 10'b1000010111;
    n950[29] = 10'b1000010110;
    n950[28] = 10'b1000010101;
    n950[27] = 10'b1000010101;
    n950[26] = 10'b1000010100;
    n950[25] = 10'b1000010011;
    n950[24] = 10'b1000010010;
    n950[23] = 10'b1000010010;
    n950[22] = 10'b1000010001;
    n950[21] = 10'b1000010000;
    n950[20] = 10'b1000001111;
    n950[19] = 10'b1000001110;
    n950[18] = 10'b1000001110;
    n950[17] = 10'b1000001101;
    n950[16] = 10'b1000001100;
    n950[15] = 10'b1000001011;
    n950[14] = 10'b1000001010;
    n950[13] = 10'b1000001010;
    n950[12] = 10'b1000001001;
    n950[11] = 10'b1000001000;
    n950[10] = 10'b1000000111;
    n950[9] = 10'b1000000111;
    n950[8] = 10'b1000000110;
    n950[7] = 10'b1000000101;
    n950[6] = 10'b1000000100;
    n950[5] = 10'b1000000011;
    n950[4] = 10'b1000000011;
    n950[3] = 10'b1000000010;
    n950[2] = 10'b1000000001;
    n950[1] = 10'b1000000000;
    n950[0] = 10'b1000000000;
    end
  assign n952 = n950[n921];
  /* ../../vhdl/src/phase_to_amplitude.vhd:47:28  */
endmodule

module phase_accumulator
  (input  clock_i,
   input  reset_i,
   input  [31:0] phase_increment_i,
   input  phase_sync_strobe_i,
   input  phase_set_strobe_i,
   input  [31:0] phase_value_i,
   output [31:0] phase_o);
  wire [31:0] phase_increment_reg;
  wire [31:0] phase_increment_next;
  wire [31:0] phase_reg;
  wire [31:0] phase_next;
  wire [32:0] n885;
  wire [32:0] n887;
  wire [32:0] n888;
  wire [31:0] n889;
  wire [31:0] n890;
  wire [31:0] n893;
  reg [31:0] n905;
  reg [31:0] n906;
  assign phase_o = phase_reg; //(module output)
  /* ../../vhdl/src/phase_accumulator.vhd:19:12  */
  assign phase_increment_reg = n905; // (signal)
  /* ../../vhdl/src/phase_accumulator.vhd:20:12  */
  assign phase_increment_next = phase_increment_i; // (signal)
  /* ../../vhdl/src/phase_accumulator.vhd:21:12  */
  assign phase_reg = n906; // (signal)
  /* ../../vhdl/src/phase_accumulator.vhd:22:12  */
  assign phase_next = n893; // (signal)
  /* ../../vhdl/src/phase_accumulator.vhd:39:33  */
  assign n885 = {1'b0, phase_reg};
  /* ../../vhdl/src/phase_accumulator.vhd:39:53  */
  assign n887 = {1'b0, phase_increment_reg};
  /* ../../vhdl/src/phase_accumulator.vhd:39:46  */
  assign n888 = n885 + n887;
  /* ../../vhdl/src/phase_accumulator.vhd:40:38  */
  assign n889 = n888[31:0]; // extract
  /* ../../vhdl/src/phase_accumulator.vhd:36:17  */
  assign n890 = phase_set_strobe_i ? phase_value_i : n889;
  /* ../../vhdl/src/phase_accumulator.vhd:34:17  */
  assign n893 = phase_sync_strobe_i ? 32'b00000000000000000000000000000000 : n890;
  /* ../../vhdl/src/phase_accumulator.vhd:50:17  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n905 <= 32'b00000000000000000000000000000000;
    else
      n905 <= phase_increment_next;
  /* ../../vhdl/src/phase_accumulator.vhd:50:17  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n906 <= 32'b00000000000000000000000000000000;
    else
      n906 <= phase_next;
endmodule

module sigma_delta_modulator
  (input  clock_i,
   input  reset_i,
   input  [9:0] sample_i,
   output bit_o);
  wire [9:0] stage_1_accumulator_1_reg;
  wire [9:0] stage_1_accumulator_1_next;
  wire [9:0] stage_1_accumulator_2_reg;
  wire [9:0] stage_1_accumulator_2_next;
  wire [1:0] stage_1_clock_divider_reg;
  wire [1:0] stage_1_clock_divider_next;
  wire [1:0] stage_1_output_reg;
  wire [1:0] stage_1_output_next;
  wire [1:0] stage_2_accumulator_reg;
  wire [1:0] stage_2_accumulator_next;
  wire bit_reg;
  wire bit_next;
  wire n820;
  wire [11:0] n822;
  wire [10:0] n824;
  wire [11:0] n826;
  wire [11:0] n828;
  wire [11:0] n829;
  wire [11:0] n831;
  wire [11:0] n832;
  wire [1:0] n833;
  wire [9:0] n834;
  wire [9:0] n835;
  wire [9:0] n836;
  wire [1:0] n837;
  wire [1:0] n845;
  wire [2:0] n847;
  wire [2:0] n849;
  wire [2:0] n850;
  wire n851;
  wire [1:0] n852;
  reg [9:0] n875;
  reg [9:0] n876;
  reg [1:0] n877;
  reg [1:0] n878;
  reg [1:0] n879;
  reg n880;
  assign bit_o = bit_reg; //(module output)
  /* ../../vhdl/src/sigma_delta_modulator.vhd:16:10  */
  assign stage_1_accumulator_1_reg = n875; // (signal)
  /* ../../vhdl/src/sigma_delta_modulator.vhd:17:10  */
  assign stage_1_accumulator_1_next = n835; // (signal)
  /* ../../vhdl/src/sigma_delta_modulator.vhd:18:10  */
  assign stage_1_accumulator_2_reg = n876; // (signal)
  /* ../../vhdl/src/sigma_delta_modulator.vhd:19:10  */
  assign stage_1_accumulator_2_next = n836; // (signal)
  /* ../../vhdl/src/sigma_delta_modulator.vhd:20:10  */
  assign stage_1_clock_divider_reg = n877; // (signal)
  /* ../../vhdl/src/sigma_delta_modulator.vhd:21:10  */
  assign stage_1_clock_divider_next = n845; // (signal)
  /* ../../vhdl/src/sigma_delta_modulator.vhd:22:10  */
  assign stage_1_output_reg = n878; // (signal)
  /* ../../vhdl/src/sigma_delta_modulator.vhd:23:10  */
  assign stage_1_output_next = n837; // (signal)
  /* ../../vhdl/src/sigma_delta_modulator.vhd:24:10  */
  assign stage_2_accumulator_reg = n879; // (signal)
  /* ../../vhdl/src/sigma_delta_modulator.vhd:25:10  */
  assign stage_2_accumulator_next = n852; // (signal)
  /* ../../vhdl/src/sigma_delta_modulator.vhd:26:10  */
  assign bit_reg = n880; // (signal)
  /* ../../vhdl/src/sigma_delta_modulator.vhd:27:10  */
  assign bit_next = n851; // (signal)
  /* ../../vhdl/src/sigma_delta_modulator.vhd:48:34  */
  assign n820 = stage_1_clock_divider_reg == 2'b00;
  /* ../../vhdl/src/sigma_delta_modulator.vhd:49:30  */
  assign n822 = {2'b00, sample_i};
  /* ../../vhdl/src/sigma_delta_modulator.vhd:50:41  */
  assign n824 = {1'b0, stage_1_accumulator_1_reg};
  /* ../../vhdl/src/sigma_delta_modulator.vhd:50:69  */
  assign n826 = {n824, 1'b0};
  /* ../../vhdl/src/sigma_delta_modulator.vhd:52:33  */
  assign n828 = {2'b00, stage_1_accumulator_2_reg};
  /* ../../vhdl/src/sigma_delta_modulator.vhd:53:30  */
  assign n829 = n822 + n826;
  /* ../../vhdl/src/sigma_delta_modulator.vhd:53:58  */
  assign n831 = n829 + 12'b010000000000;
  /* ../../vhdl/src/sigma_delta_modulator.vhd:53:73  */
  assign n832 = n831 - n828;
  /* ../../vhdl/src/sigma_delta_modulator.vhd:55:35  */
  assign n833 = n832[11:10]; // extract
  /* ../../vhdl/src/sigma_delta_modulator.vhd:56:42  */
  assign n834 = n832[9:0]; // extract
  /* ../../vhdl/src/sigma_delta_modulator.vhd:48:5  */
  assign n835 = n820 ? n834 : stage_1_accumulator_1_reg;
  /* ../../vhdl/src/sigma_delta_modulator.vhd:48:5  */
  assign n836 = n820 ? stage_1_accumulator_1_reg : stage_1_accumulator_2_reg;
  /* ../../vhdl/src/sigma_delta_modulator.vhd:48:5  */
  assign n837 = n820 ? n833 : stage_1_output_reg;
  /* ../../vhdl/src/sigma_delta_modulator.vhd:60:61  */
  assign n845 = stage_1_clock_divider_reg + 2'b01;
  /* ../../vhdl/src/sigma_delta_modulator.vhd:61:19  */
  assign n847 = {1'b0, stage_2_accumulator_reg};
  /* ../../vhdl/src/sigma_delta_modulator.vhd:61:53  */
  assign n849 = {1'b0, stage_1_output_reg};
  /* ../../vhdl/src/sigma_delta_modulator.vhd:61:46  */
  assign n850 = n847 + n849;
  /* ../../vhdl/src/sigma_delta_modulator.vhd:62:22  */
  assign n851 = n850[2]; // extract
  /* ../../vhdl/src/sigma_delta_modulator.vhd:63:39  */
  assign n852 = n850[1:0]; // extract
  /* ../../vhdl/src/sigma_delta_modulator.vhd:75:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n875 <= 10'b0000000000;
    else
      n875 <= stage_1_accumulator_1_next;
  /* ../../vhdl/src/sigma_delta_modulator.vhd:75:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n876 <= 10'b0000000000;
    else
      n876 <= stage_1_accumulator_2_next;
  /* ../../vhdl/src/sigma_delta_modulator.vhd:75:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n877 <= 2'b00;
    else
      n877 <= stage_1_clock_divider_next;
  /* ../../vhdl/src/sigma_delta_modulator.vhd:75:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n878 <= 2'b00;
    else
      n878 <= stage_1_output_next;
  /* ../../vhdl/src/sigma_delta_modulator.vhd:75:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n879 <= 2'b00;
    else
      n879 <= stage_2_accumulator_next;
  /* ../../vhdl/src/sigma_delta_modulator.vhd:75:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n880 <= 1'b0;
    else
      n880 <= bit_next;
endmodule

module direct_digital_synthesis
  (input  clock_i,
   input  reset_i,
   input  [31:0] phase_increment_i,
   input  phase_sync_strobe_i,
   input  phase_set_strobe_i,
   input  [31:0] phase_value_i,
   output [9:0] sample_o);
  wire [31:0] phase;
  wire [9:0] \phase_to_amplitude_instance.amplitude_o ;
  assign sample_o = \phase_to_amplitude_instance.amplitude_o ; //(module output)
  /* ../../vhdl/src/direct_digital_synthesis.vhd:24:5  */
  phase_accumulator phase_accumulator_instance (
    .clock_i(clock_i),
    .reset_i(reset_i),
    .phase_increment_i(phase_increment_i),
    .phase_sync_strobe_i(phase_sync_strobe_i),
    .phase_set_strobe_i(phase_set_strobe_i),
    .phase_value_i(phase_value_i),
    .phase_o(phase));
  /* ../../vhdl/src/direct_digital_synthesis.vhd:35:5  */
  phase_to_amplitude phase_to_amplitude_instance (
    .clock_i(clock_i),
    .reset_i(reset_i),
    .phase_i(phase),
    .amplitude_o(\phase_to_amplitude_instance.amplitude_o ));
endmodule

module channel
  (input  clock_i,
   input  reset_i,
   input  [31:0] phase_increment_i,
   input  phase_sync_strobe_i,
   input  phase_set_strobe_i,
   input  [31:0] phase_value_i,
   output wave_o);
  wire [9:0] sample;
  wire \sigma_delta_modulator_instance.bit_o ;
  assign wave_o = \sigma_delta_modulator_instance.bit_o ; //(module output)
  /* ../../vhdl/src/channel.vhd:22:5  */
  direct_digital_synthesis direct_digital_synthesis_instance (
    .clock_i(clock_i),
    .reset_i(reset_i),
    .phase_increment_i(phase_increment_i),
    .phase_sync_strobe_i(phase_sync_strobe_i),
    .phase_set_strobe_i(phase_set_strobe_i),
    .phase_value_i(phase_value_i),
    .sample_o(sample));
  /* ../../vhdl/src/channel.vhd:33:6  */
  sigma_delta_modulator sigma_delta_modulator_instance (
    .clock_i(clock_i),
    .reset_i(reset_i),
    .sample_i(sample),
    .bit_o(\sigma_delta_modulator_instance.bit_o ));
endmodule

module uart_tx
  (input  clock_i,
   input  reset_i,
   input  tx_data_valid_i,
   input  [7:0] tx_data_i,
   output tx_active_o,
   output serial_o,
   output tx_done_o);
  wire [1:0] state_reg;
  wire [1:0] state_next;
  wire [8:0] bit_clock_counter_reg;
  wire [8:0] bit_clock_counter_next;
  wire [2:0] bit_index_reg;
  wire [2:0] bit_index_next;
  wire [7:0] tx_shift_reg;
  wire [7:0] tx_shift_next;
  wire tx_done_reg;
  wire tx_done_next;
  wire tx_active_reg;
  wire tx_active_next;
  wire serial_out_reg;
  wire serial_out_next;
  wire [1:0] n676;
  wire [8:0] n679;
  wire [7:0] n681;
  wire n684;
  wire n687;
  wire [31:0] n688;
  wire n690;
  wire [31:0] n691;
  wire [31:0] n693;
  wire [8:0] n694;
  wire [1:0] n696;
  wire [8:0] n698;
  wire n700;
  wire n701;
  wire [31:0] n702;
  wire n704;
  wire [6:0] n705;
  wire [7:0] n707;
  wire [31:0] n708;
  wire n710;
  wire [31:0] n711;
  wire [31:0] n713;
  wire [2:0] n714;
  wire [1:0] n716;
  wire [2:0] n718;
  wire [31:0] n719;
  wire [31:0] n721;
  wire [8:0] n722;
  wire [1:0] n723;
  wire [8:0] n725;
  wire [2:0] n726;
  wire [7:0] n727;
  wire n729;
  wire [31:0] n730;
  wire n732;
  wire [31:0] n733;
  wire [31:0] n735;
  wire [8:0] n736;
  wire [1:0] n738;
  wire [8:0] n739;
  wire n742;
  wire n745;
  wire n748;
  wire [3:0] n749;
  reg [1:0] n751;
  reg [8:0] n753;
  reg [2:0] n756;
  reg [7:0] n758;
  reg n761;
  reg n766;
  reg n771;
  reg [1:0] n797;
  reg [8:0] n798;
  reg [2:0] n799;
  reg [7:0] n800;
  reg n801;
  reg n802;
  reg n803;
  assign tx_active_o = tx_active_reg; //(module output)
  assign serial_o = serial_out_reg; //(module output)
  assign tx_done_o = tx_done_reg; //(module output)
  /* ../../vhdl/src/UART_TX.vhd:20:10  */
  assign state_reg = n797; // (signal)
  /* ../../vhdl/src/UART_TX.vhd:21:10  */
  assign state_next = n751; // (signal)
  /* ../../vhdl/src/UART_TX.vhd:22:10  */
  assign bit_clock_counter_reg = n798; // (signal)
  /* ../../vhdl/src/UART_TX.vhd:23:10  */
  assign bit_clock_counter_next = n753; // (signal)
  /* ../../vhdl/src/UART_TX.vhd:24:10  */
  assign bit_index_reg = n799; // (signal)
  /* ../../vhdl/src/UART_TX.vhd:25:10  */
  assign bit_index_next = n756; // (signal)
  /* ../../vhdl/src/UART_TX.vhd:26:10  */
  assign tx_shift_reg = n800; // (signal)
  /* ../../vhdl/src/UART_TX.vhd:27:10  */
  assign tx_shift_next = n758; // (signal)
  /* ../../vhdl/src/UART_TX.vhd:28:10  */
  assign tx_done_reg = n801; // (signal)
  /* ../../vhdl/src/UART_TX.vhd:29:10  */
  assign tx_done_next = n761; // (signal)
  /* ../../vhdl/src/UART_TX.vhd:30:10  */
  assign tx_active_reg = n802; // (signal)
  /* ../../vhdl/src/UART_TX.vhd:31:10  */
  assign tx_active_next = n766; // (signal)
  /* ../../vhdl/src/UART_TX.vhd:32:10  */
  assign serial_out_reg = n803; // (signal)
  /* ../../vhdl/src/UART_TX.vhd:33:10  */
  assign serial_out_next = n771; // (signal)
  /* ../../vhdl/src/UART_TX.vhd:54:9  */
  assign n676 = tx_data_valid_i ? 2'b01 : state_reg;
  /* ../../vhdl/src/UART_TX.vhd:54:9  */
  assign n679 = tx_data_valid_i ? 9'b100010101 : 9'b000000000;
  /* ../../vhdl/src/UART_TX.vhd:54:9  */
  assign n681 = tx_data_valid_i ? tx_data_i : tx_shift_reg;
  /* ../../vhdl/src/UART_TX.vhd:54:9  */
  assign n684 = tx_data_valid_i ? 1'b1 : 1'b0;
  /* ../../vhdl/src/UART_TX.vhd:49:7  */
  assign n687 = state_reg == 2'b00;
  /* ../../vhdl/src/UART_TX.vhd:64:34  */
  assign n688 = {23'b0, bit_clock_counter_reg};  //  uext
  /* ../../vhdl/src/UART_TX.vhd:64:34  */
  assign n690 = n688 == 32'b00000000000000000000000000000000;
  /* ../../vhdl/src/UART_TX.vhd:68:59  */
  assign n691 = {23'b0, bit_clock_counter_reg};  //  uext
  /* ../../vhdl/src/UART_TX.vhd:68:59  */
  assign n693 = n691 - 32'b00000000000000000000000000000001;
  /* ../../vhdl/src/UART_TX.vhd:68:37  */
  assign n694 = n693[8:0];  // trunc
  /* ../../vhdl/src/UART_TX.vhd:64:9  */
  assign n696 = n690 ? 2'b10 : state_reg;
  /* ../../vhdl/src/UART_TX.vhd:64:9  */
  assign n698 = n690 ? 9'b100010101 : n694;
  /* ../../vhdl/src/UART_TX.vhd:61:7  */
  assign n700 = state_reg == 2'b01;
  /* ../../vhdl/src/UART_TX.vhd:73:40  */
  assign n701 = tx_shift_reg[0]; // extract
  /* ../../vhdl/src/UART_TX.vhd:74:34  */
  assign n702 = {23'b0, bit_clock_counter_reg};  //  uext
  /* ../../vhdl/src/UART_TX.vhd:74:34  */
  assign n704 = n702 == 32'b00000000000000000000000000000000;
  /* ../../vhdl/src/UART_TX.vhd:76:46  */
  assign n705 = tx_shift_reg[7:1]; // extract
  /* ../../vhdl/src/UART_TX.vhd:76:32  */
  assign n707 = {1'b0, n705};
  /* ../../vhdl/src/UART_TX.vhd:77:28  */
  assign n708 = {29'b0, bit_index_reg};  //  uext
  /* ../../vhdl/src/UART_TX.vhd:77:28  */
  assign n710 = $signed(n708) < $signed(32'b00000000000000000000000000000111);
  /* ../../vhdl/src/UART_TX.vhd:78:45  */
  assign n711 = {29'b0, bit_index_reg};  //  uext
  /* ../../vhdl/src/UART_TX.vhd:78:45  */
  assign n713 = n711 + 32'b00000000000000000000000000000001;
  /* ../../vhdl/src/UART_TX.vhd:78:31  */
  assign n714 = n713[2:0];  // trunc
  /* ../../vhdl/src/UART_TX.vhd:77:11  */
  assign n716 = n710 ? state_reg : 2'b11;
  /* ../../vhdl/src/UART_TX.vhd:77:11  */
  assign n718 = n710 ? n714 : 3'b000;
  /* ../../vhdl/src/UART_TX.vhd:84:59  */
  assign n719 = {23'b0, bit_clock_counter_reg};  //  uext
  /* ../../vhdl/src/UART_TX.vhd:84:59  */
  assign n721 = n719 - 32'b00000000000000000000000000000001;
  /* ../../vhdl/src/UART_TX.vhd:84:37  */
  assign n722 = n721[8:0];  // trunc
  /* ../../vhdl/src/UART_TX.vhd:74:9  */
  assign n723 = n704 ? n716 : state_reg;
  /* ../../vhdl/src/UART_TX.vhd:74:9  */
  assign n725 = n704 ? 9'b100010101 : n722;
  /* ../../vhdl/src/UART_TX.vhd:74:9  */
  assign n726 = n704 ? n718 : bit_index_reg;
  /* ../../vhdl/src/UART_TX.vhd:74:9  */
  assign n727 = n704 ? n707 : tx_shift_reg;
  /* ../../vhdl/src/UART_TX.vhd:71:7  */
  assign n729 = state_reg == 2'b10;
  /* ../../vhdl/src/UART_TX.vhd:90:34  */
  assign n730 = {23'b0, bit_clock_counter_reg};  //  uext
  /* ../../vhdl/src/UART_TX.vhd:90:34  */
  assign n732 = n730 == 32'b00000000000000000000000000000000;
  /* ../../vhdl/src/UART_TX.vhd:95:59  */
  assign n733 = {23'b0, bit_clock_counter_reg};  //  uext
  /* ../../vhdl/src/UART_TX.vhd:95:59  */
  assign n735 = n733 - 32'b00000000000000000000000000000001;
  /* ../../vhdl/src/UART_TX.vhd:95:37  */
  assign n736 = n735[8:0];  // trunc
  /* ../../vhdl/src/UART_TX.vhd:90:9  */
  assign n738 = n732 ? 2'b00 : state_reg;
  /* ../../vhdl/src/UART_TX.vhd:90:9  */
  assign n739 = n732 ? bit_clock_counter_reg : n736;
  /* ../../vhdl/src/UART_TX.vhd:90:9  */
  assign n742 = n732 ? 1'b1 : 1'b0;
  /* ../../vhdl/src/UART_TX.vhd:90:9  */
  assign n745 = n732 ? 1'b0 : 1'b1;
  /* ../../vhdl/src/UART_TX.vhd:87:7  */
  assign n748 = state_reg == 2'b11;
  assign n749 = {n748, n729, n700, n687};
  /* ../../vhdl/src/UART_TX.vhd:47:5  */
  always @*
    case (n749)
      4'b1000: n751 = n738;
      4'b0100: n751 = n723;
      4'b0010: n751 = n696;
      4'b0001: n751 = n676;
      default: n751 = 2'b00;
    endcase
  /* ../../vhdl/src/UART_TX.vhd:47:5  */
  always @*
    case (n749)
      4'b1000: n753 = n739;
      4'b0100: n753 = n725;
      4'b0010: n753 = n698;
      4'b0001: n753 = n679;
      default: n753 = 9'b000000000;
    endcase
  /* ../../vhdl/src/UART_TX.vhd:47:5  */
  always @*
    case (n749)
      4'b1000: n756 = bit_index_reg;
      4'b0100: n756 = n726;
      4'b0010: n756 = bit_index_reg;
      4'b0001: n756 = 3'b000;
      default: n756 = 3'b000;
    endcase
  /* ../../vhdl/src/UART_TX.vhd:47:5  */
  always @*
    case (n749)
      4'b1000: n758 = tx_shift_reg;
      4'b0100: n758 = n727;
      4'b0010: n758 = tx_shift_reg;
      4'b0001: n758 = n681;
      default: n758 = 8'b00000000;
    endcase
  /* ../../vhdl/src/UART_TX.vhd:47:5  */
  always @*
    case (n749)
      4'b1000: n761 = n742;
      4'b0100: n761 = 1'b0;
      4'b0010: n761 = 1'b0;
      4'b0001: n761 = 1'b0;
      default: n761 = 1'b0;
    endcase
  /* ../../vhdl/src/UART_TX.vhd:47:5  */
  always @*
    case (n749)
      4'b1000: n766 = n745;
      4'b0100: n766 = 1'b1;
      4'b0010: n766 = 1'b1;
      4'b0001: n766 = n684;
      default: n766 = 1'b0;
    endcase
  /* ../../vhdl/src/UART_TX.vhd:47:5  */
  always @*
    case (n749)
      4'b1000: n771 = 1'b1;
      4'b0100: n771 = n701;
      4'b0010: n771 = 1'b0;
      4'b0001: n771 = 1'b1;
      default: n771 = 1'b1;
    endcase
  /* ../../vhdl/src/UART_TX.vhd:119:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n797 <= 2'b00;
    else
      n797 <= state_next;
  /* ../../vhdl/src/UART_TX.vhd:119:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n798 <= 9'b000000000;
    else
      n798 <= bit_clock_counter_next;
  /* ../../vhdl/src/UART_TX.vhd:119:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n799 <= 3'b000;
    else
      n799 <= bit_index_next;
  /* ../../vhdl/src/UART_TX.vhd:119:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n800 <= 8'b00000000;
    else
      n800 <= tx_shift_next;
  /* ../../vhdl/src/UART_TX.vhd:119:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n801 <= 1'b0;
    else
      n801 <= tx_done_next;
  /* ../../vhdl/src/UART_TX.vhd:119:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n802 <= 1'b0;
    else
      n802 <= tx_active_next;
  /* ../../vhdl/src/UART_TX.vhd:119:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n803 <= 1'b1;
    else
      n803 <= serial_out_next;
endmodule

module uart_rx
  (input  clock_i,
   input  reset_i,
   input  serial_i,
   output data_valid_o,
   output [7:0] rx_byte_o);
  wire [1:0] state_reg;
  wire [1:0] state_next;
  wire [8:0] bit_clock_counter_reg;
  wire [8:0] bit_clock_counter_next;
  wire [2:0] bit_index_reg;
  wire [2:0] bit_index_next;
  wire [7:0] rx_shift_reg;
  wire [7:0] rx_shift_next;
  wire data_valid_reg;
  wire data_valid_next;
  wire [7:0] rx_output_reg;
  wire [7:0] rx_output_next;
  wire serial_sync1_reg;
  wire serial_sync1_next;
  wire serial_sync2_reg;
  wire serial_sync2_next;
  wire n546;
  wire [1:0] n549;
  wire [8:0] n552;
  wire n555;
  wire [31:0] n556;
  wire n558;
  wire n559;
  wire [1:0] n562;
  wire [8:0] n564;
  wire [31:0] n565;
  wire [31:0] n567;
  wire [8:0] n568;
  wire [1:0] n569;
  wire [8:0] n570;
  wire n572;
  wire [31:0] n573;
  wire n575;
  wire [6:0] n576;
  wire [7:0] n577;
  wire [31:0] n578;
  wire n580;
  wire [31:0] n581;
  wire [31:0] n583;
  wire [2:0] n584;
  wire [1:0] n587;
  wire [2:0] n589;
  wire [31:0] n590;
  wire [31:0] n592;
  wire [8:0] n593;
  wire [1:0] n594;
  wire [8:0] n596;
  wire [2:0] n597;
  wire [7:0] n598;
  wire n600;
  wire [31:0] n601;
  wire n603;
  wire n606;
  wire [7:0] n607;
  wire [31:0] n608;
  wire [31:0] n610;
  wire [8:0] n611;
  wire [1:0] n613;
  wire [8:0] n614;
  wire n616;
  wire n617;
  wire n619;
  wire [3:0] n620;
  reg [1:0] n622;
  reg [8:0] n624;
  reg [2:0] n627;
  reg [7:0] n629;
  reg n632;
  reg [7:0] n634;
  reg [1:0] n663;
  reg [8:0] n664;
  reg [2:0] n665;
  reg [7:0] n666;
  reg n667;
  reg [7:0] n668;
  reg n669;
  reg n670;
  assign data_valid_o = data_valid_reg; //(module output)
  assign rx_byte_o = rx_output_reg; //(module output)
  /* ../../vhdl/src/UART_RX.vhd:18:10  */
  assign state_reg = n663; // (signal)
  /* ../../vhdl/src/UART_RX.vhd:19:10  */
  assign state_next = n622; // (signal)
  /* ../../vhdl/src/UART_RX.vhd:20:10  */
  assign bit_clock_counter_reg = n664; // (signal)
  /* ../../vhdl/src/UART_RX.vhd:21:10  */
  assign bit_clock_counter_next = n624; // (signal)
  /* ../../vhdl/src/UART_RX.vhd:22:10  */
  assign bit_index_reg = n665; // (signal)
  /* ../../vhdl/src/UART_RX.vhd:23:10  */
  assign bit_index_next = n627; // (signal)
  /* ../../vhdl/src/UART_RX.vhd:24:10  */
  assign rx_shift_reg = n666; // (signal)
  /* ../../vhdl/src/UART_RX.vhd:25:10  */
  assign rx_shift_next = n629; // (signal)
  /* ../../vhdl/src/UART_RX.vhd:26:10  */
  assign data_valid_reg = n667; // (signal)
  /* ../../vhdl/src/UART_RX.vhd:27:10  */
  assign data_valid_next = n632; // (signal)
  /* ../../vhdl/src/UART_RX.vhd:28:10  */
  assign rx_output_reg = n668; // (signal)
  /* ../../vhdl/src/UART_RX.vhd:29:10  */
  assign rx_output_next = n634; // (signal)
  /* ../../vhdl/src/UART_RX.vhd:30:10  */
  assign serial_sync1_reg = n669; // (signal)
  /* ../../vhdl/src/UART_RX.vhd:31:10  */
  assign serial_sync1_next = serial_i; // (signal)
  /* ../../vhdl/src/UART_RX.vhd:32:10  */
  assign serial_sync2_reg = n670; // (signal)
  /* ../../vhdl/src/UART_RX.vhd:33:10  */
  assign serial_sync2_next = serial_sync1_reg; // (signal)
  /* ../../vhdl/src/UART_RX.vhd:56:29  */
  assign n546 = ~serial_sync2_reg;
  /* ../../vhdl/src/UART_RX.vhd:56:9  */
  assign n549 = n546 ? 2'b01 : 2'b00;
  /* ../../vhdl/src/UART_RX.vhd:56:9  */
  assign n552 = n546 ? 9'b010001010 : 9'b000000000;
  /* ../../vhdl/src/UART_RX.vhd:53:7  */
  assign n555 = state_reg == 2'b00;
  /* ../../vhdl/src/UART_RX.vhd:64:34  */
  assign n556 = {23'b0, bit_clock_counter_reg};  //  uext
  /* ../../vhdl/src/UART_RX.vhd:64:34  */
  assign n558 = n556 == 32'b00000000000000000000000000000000;
  /* ../../vhdl/src/UART_RX.vhd:65:32  */
  assign n559 = ~serial_sync2_reg;
  /* ../../vhdl/src/UART_RX.vhd:65:12  */
  assign n562 = n559 ? 2'b10 : 2'b00;
  /* ../../vhdl/src/UART_RX.vhd:65:12  */
  assign n564 = n559 ? 9'b100010101 : bit_clock_counter_reg;
  /* ../../vhdl/src/UART_RX.vhd:72:60  */
  assign n565 = {23'b0, bit_clock_counter_reg};  //  uext
  /* ../../vhdl/src/UART_RX.vhd:72:60  */
  assign n567 = n565 - 32'b00000000000000000000000000000001;
  /* ../../vhdl/src/UART_RX.vhd:72:38  */
  assign n568 = n567[8:0];  // trunc
  /* ../../vhdl/src/UART_RX.vhd:64:9  */
  assign n569 = n558 ? n562 : state_reg;
  /* ../../vhdl/src/UART_RX.vhd:64:9  */
  assign n570 = n558 ? n564 : n568;
  /* ../../vhdl/src/UART_RX.vhd:63:7  */
  assign n572 = state_reg == 2'b01;
  /* ../../vhdl/src/UART_RX.vhd:76:34  */
  assign n573 = {23'b0, bit_clock_counter_reg};  //  uext
  /* ../../vhdl/src/UART_RX.vhd:76:34  */
  assign n575 = n573 == 32'b00000000000000000000000000000000;
  /* ../../vhdl/src/UART_RX.vhd:78:59  */
  assign n576 = rx_shift_reg[7:1]; // extract
  /* ../../vhdl/src/UART_RX.vhd:78:45  */
  assign n577 = {serial_sync2_reg, n576};
  /* ../../vhdl/src/UART_RX.vhd:79:28  */
  assign n578 = {29'b0, bit_index_reg};  //  uext
  /* ../../vhdl/src/UART_RX.vhd:79:28  */
  assign n580 = $signed(n578) < $signed(32'b00000000000000000000000000000111);
  /* ../../vhdl/src/UART_RX.vhd:80:45  */
  assign n581 = {29'b0, bit_index_reg};  //  uext
  /* ../../vhdl/src/UART_RX.vhd:80:45  */
  assign n583 = n581 + 32'b00000000000000000000000000000001;
  /* ../../vhdl/src/UART_RX.vhd:80:31  */
  assign n584 = n583[2:0];  // trunc
  /* ../../vhdl/src/UART_RX.vhd:79:11  */
  assign n587 = n580 ? 2'b10 : 2'b11;
  /* ../../vhdl/src/UART_RX.vhd:79:11  */
  assign n589 = n580 ? n584 : 3'b000;
  /* ../../vhdl/src/UART_RX.vhd:87:59  */
  assign n590 = {23'b0, bit_clock_counter_reg};  //  uext
  /* ../../vhdl/src/UART_RX.vhd:87:59  */
  assign n592 = n590 - 32'b00000000000000000000000000000001;
  /* ../../vhdl/src/UART_RX.vhd:87:37  */
  assign n593 = n592[8:0];  // trunc
  /* ../../vhdl/src/UART_RX.vhd:76:9  */
  assign n594 = n575 ? n587 : state_reg;
  /* ../../vhdl/src/UART_RX.vhd:76:9  */
  assign n596 = n575 ? 9'b100010101 : n593;
  /* ../../vhdl/src/UART_RX.vhd:76:9  */
  assign n597 = n575 ? n589 : bit_index_reg;
  /* ../../vhdl/src/UART_RX.vhd:76:9  */
  assign n598 = n575 ? n577 : rx_shift_reg;
  /* ../../vhdl/src/UART_RX.vhd:75:7  */
  assign n600 = state_reg == 2'b10;
  /* ../../vhdl/src/UART_RX.vhd:91:34  */
  assign n601 = {23'b0, bit_clock_counter_reg};  //  uext
  /* ../../vhdl/src/UART_RX.vhd:91:34  */
  assign n603 = n601 == 32'b00000000000000000000000000000000;
  /* ../../vhdl/src/UART_RX.vhd:92:11  */
  assign n606 = serial_sync2_reg ? 1'b1 : 1'b0;
  /* ../../vhdl/src/UART_RX.vhd:91:9  */
  assign n607 = n617 ? rx_shift_reg : rx_output_reg;
  /* ../../vhdl/src/UART_RX.vhd:98:59  */
  assign n608 = {23'b0, bit_clock_counter_reg};  //  uext
  /* ../../vhdl/src/UART_RX.vhd:98:59  */
  assign n610 = n608 - 32'b00000000000000000000000000000001;
  /* ../../vhdl/src/UART_RX.vhd:98:37  */
  assign n611 = n610[8:0];  // trunc
  /* ../../vhdl/src/UART_RX.vhd:91:9  */
  assign n613 = n603 ? 2'b00 : state_reg;
  /* ../../vhdl/src/UART_RX.vhd:91:9  */
  assign n614 = n603 ? bit_clock_counter_reg : n611;
  /* ../../vhdl/src/UART_RX.vhd:91:9  */
  assign n616 = n603 ? n606 : 1'b0;
  /* ../../vhdl/src/UART_RX.vhd:91:9  */
  assign n617 = serial_sync2_reg & n603;
  /* ../../vhdl/src/UART_RX.vhd:90:7  */
  assign n619 = state_reg == 2'b11;
  assign n620 = {n619, n600, n572, n555};
  /* ../../vhdl/src/UART_RX.vhd:51:5  */
  always @*
    case (n620)
      4'b1000: n622 = n613;
      4'b0100: n622 = n594;
      4'b0010: n622 = n569;
      4'b0001: n622 = n549;
      default: n622 = 2'b00;
    endcase
  /* ../../vhdl/src/UART_RX.vhd:51:5  */
  always @*
    case (n620)
      4'b1000: n624 = n614;
      4'b0100: n624 = n596;
      4'b0010: n624 = n570;
      4'b0001: n624 = n552;
      default: n624 = 9'b000000000;
    endcase
  /* ../../vhdl/src/UART_RX.vhd:51:5  */
  always @*
    case (n620)
      4'b1000: n627 = bit_index_reg;
      4'b0100: n627 = n597;
      4'b0010: n627 = bit_index_reg;
      4'b0001: n627 = 3'b000;
      default: n627 = 3'b000;
    endcase
  /* ../../vhdl/src/UART_RX.vhd:51:5  */
  always @*
    case (n620)
      4'b1000: n629 = rx_shift_reg;
      4'b0100: n629 = n598;
      4'b0010: n629 = rx_shift_reg;
      4'b0001: n629 = rx_shift_reg;
      default: n629 = 8'b00000000;
    endcase
  /* ../../vhdl/src/UART_RX.vhd:51:5  */
  always @*
    case (n620)
      4'b1000: n632 = n616;
      4'b0100: n632 = 1'b0;
      4'b0010: n632 = 1'b0;
      4'b0001: n632 = 1'b0;
      default: n632 = 1'b0;
    endcase
  /* ../../vhdl/src/UART_RX.vhd:51:5  */
  always @*
    case (n620)
      4'b1000: n634 = n607;
      4'b0100: n634 = rx_output_reg;
      4'b0010: n634 = rx_output_reg;
      4'b0001: n634 = rx_output_reg;
      default: n634 = rx_output_reg;
    endcase
  /* ../../vhdl/src/UART_RX.vhd:121:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n663 <= 2'b00;
    else
      n663 <= state_next;
  /* ../../vhdl/src/UART_RX.vhd:121:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n664 <= 9'b000000000;
    else
      n664 <= bit_clock_counter_next;
  /* ../../vhdl/src/UART_RX.vhd:121:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n665 <= 3'b000;
    else
      n665 <= bit_index_next;
  /* ../../vhdl/src/UART_RX.vhd:121:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n666 <= 8'b00000000;
    else
      n666 <= rx_shift_next;
  /* ../../vhdl/src/UART_RX.vhd:121:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n667 <= 1'b0;
    else
      n667 <= data_valid_next;
  /* ../../vhdl/src/UART_RX.vhd:121:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n668 <= 8'b00000000;
    else
      n668 <= rx_output_next;
  /* ../../vhdl/src/UART_RX.vhd:121:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n669 <= 1'b1;
    else
      n669 <= serial_sync1_next;
  /* ../../vhdl/src/UART_RX.vhd:121:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n670 <= 1'b1;
    else
      n670 <= serial_sync2_next;
endmodule

module synthesizer
  (input  clock_i,
   input  reset_i,
   input  [255:0] phase_increment_i,
   input  [255:0] phase_value_i,
   input  [7:0] phase_sync_strobe_i,
   input  [7:0] phase_set_strobe_i,
   output [7:0] waves_o);
  wire \gen_channels_n1_channel_inst.wave_o ;
  wire [31:0] n502;
  wire n503;
  wire n504;
  wire [31:0] n505;
  wire \gen_channels_n2_channel_inst.wave_o ;
  wire [31:0] n507;
  wire n508;
  wire n509;
  wire [31:0] n510;
  wire \gen_channels_n3_channel_inst.wave_o ;
  wire [31:0] n512;
  wire n513;
  wire n514;
  wire [31:0] n515;
  wire \gen_channels_n4_channel_inst.wave_o ;
  wire [31:0] n517;
  wire n518;
  wire n519;
  wire [31:0] n520;
  wire \gen_channels_n5_channel_inst.wave_o ;
  wire [31:0] n522;
  wire n523;
  wire n524;
  wire [31:0] n525;
  wire \gen_channels_n6_channel_inst.wave_o ;
  wire [31:0] n527;
  wire n528;
  wire n529;
  wire [31:0] n530;
  wire \gen_channels_n7_channel_inst.wave_o ;
  wire [31:0] n532;
  wire n533;
  wire n534;
  wire [31:0] n535;
  wire \gen_channels_n8_channel_inst.wave_o ;
  wire [31:0] n537;
  wire n538;
  wire n539;
  wire [31:0] n540;
  wire [7:0] n542;
  assign waves_o = n542; //(module output)
  /* ../../vhdl/src/synthesizer.vhd:21:9  */
  channel gen_channels_n1_channel_inst (
    .clock_i(clock_i),
    .reset_i(reset_i),
    .phase_increment_i(n502),
    .phase_sync_strobe_i(n503),
    .phase_set_strobe_i(n504),
    .phase_value_i(n505),
    .wave_o(\gen_channels_n1_channel_inst.wave_o ));
  /* ../../vhdl/src/synthesizer.vhd:25:55  */
  assign n502 = phase_increment_i[255:224]; // extract
  /* ../../vhdl/src/synthesizer.vhd:26:59  */
  assign n503 = phase_sync_strobe_i[0]; // extract
  /* ../../vhdl/src/synthesizer.vhd:27:57  */
  assign n504 = phase_set_strobe_i[0]; // extract
  /* ../../vhdl/src/synthesizer.vhd:28:47  */
  assign n505 = phase_value_i[255:224]; // extract
  /* ../../vhdl/src/synthesizer.vhd:21:9  */
  channel gen_channels_n2_channel_inst (
    .clock_i(clock_i),
    .reset_i(reset_i),
    .phase_increment_i(n507),
    .phase_sync_strobe_i(n508),
    .phase_set_strobe_i(n509),
    .phase_value_i(n510),
    .wave_o(\gen_channels_n2_channel_inst.wave_o ));
  /* ../../vhdl/src/synthesizer.vhd:25:55  */
  assign n507 = phase_increment_i[223:192]; // extract
  /* ../../vhdl/src/synthesizer.vhd:26:59  */
  assign n508 = phase_sync_strobe_i[1]; // extract
  /* ../../vhdl/src/synthesizer.vhd:27:57  */
  assign n509 = phase_set_strobe_i[1]; // extract
  /* ../../vhdl/src/synthesizer.vhd:28:47  */
  assign n510 = phase_value_i[223:192]; // extract
  /* ../../vhdl/src/synthesizer.vhd:21:9  */
  channel gen_channels_n3_channel_inst (
    .clock_i(clock_i),
    .reset_i(reset_i),
    .phase_increment_i(n512),
    .phase_sync_strobe_i(n513),
    .phase_set_strobe_i(n514),
    .phase_value_i(n515),
    .wave_o(\gen_channels_n3_channel_inst.wave_o ));
  /* ../../vhdl/src/synthesizer.vhd:25:55  */
  assign n512 = phase_increment_i[191:160]; // extract
  /* ../../vhdl/src/synthesizer.vhd:26:59  */
  assign n513 = phase_sync_strobe_i[2]; // extract
  /* ../../vhdl/src/synthesizer.vhd:27:57  */
  assign n514 = phase_set_strobe_i[2]; // extract
  /* ../../vhdl/src/synthesizer.vhd:28:47  */
  assign n515 = phase_value_i[191:160]; // extract
  /* ../../vhdl/src/synthesizer.vhd:21:9  */
  channel gen_channels_n4_channel_inst (
    .clock_i(clock_i),
    .reset_i(reset_i),
    .phase_increment_i(n517),
    .phase_sync_strobe_i(n518),
    .phase_set_strobe_i(n519),
    .phase_value_i(n520),
    .wave_o(\gen_channels_n4_channel_inst.wave_o ));
  /* ../../vhdl/src/synthesizer.vhd:25:55  */
  assign n517 = phase_increment_i[159:128]; // extract
  /* ../../vhdl/src/synthesizer.vhd:26:59  */
  assign n518 = phase_sync_strobe_i[3]; // extract
  /* ../../vhdl/src/synthesizer.vhd:27:57  */
  assign n519 = phase_set_strobe_i[3]; // extract
  /* ../../vhdl/src/synthesizer.vhd:28:47  */
  assign n520 = phase_value_i[159:128]; // extract
  /* ../../vhdl/src/synthesizer.vhd:21:9  */
  channel gen_channels_n5_channel_inst (
    .clock_i(clock_i),
    .reset_i(reset_i),
    .phase_increment_i(n522),
    .phase_sync_strobe_i(n523),
    .phase_set_strobe_i(n524),
    .phase_value_i(n525),
    .wave_o(\gen_channels_n5_channel_inst.wave_o ));
  /* ../../vhdl/src/synthesizer.vhd:25:55  */
  assign n522 = phase_increment_i[127:96]; // extract
  /* ../../vhdl/src/synthesizer.vhd:26:59  */
  assign n523 = phase_sync_strobe_i[4]; // extract
  /* ../../vhdl/src/synthesizer.vhd:27:57  */
  assign n524 = phase_set_strobe_i[4]; // extract
  /* ../../vhdl/src/synthesizer.vhd:28:47  */
  assign n525 = phase_value_i[127:96]; // extract
  /* ../../vhdl/src/synthesizer.vhd:21:9  */
  channel gen_channels_n6_channel_inst (
    .clock_i(clock_i),
    .reset_i(reset_i),
    .phase_increment_i(n527),
    .phase_sync_strobe_i(n528),
    .phase_set_strobe_i(n529),
    .phase_value_i(n530),
    .wave_o(\gen_channels_n6_channel_inst.wave_o ));
  /* ../../vhdl/src/synthesizer.vhd:25:55  */
  assign n527 = phase_increment_i[95:64]; // extract
  /* ../../vhdl/src/synthesizer.vhd:26:59  */
  assign n528 = phase_sync_strobe_i[5]; // extract
  /* ../../vhdl/src/synthesizer.vhd:27:57  */
  assign n529 = phase_set_strobe_i[5]; // extract
  /* ../../vhdl/src/synthesizer.vhd:28:47  */
  assign n530 = phase_value_i[95:64]; // extract
  /* ../../vhdl/src/synthesizer.vhd:21:9  */
  channel gen_channels_n7_channel_inst (
    .clock_i(clock_i),
    .reset_i(reset_i),
    .phase_increment_i(n532),
    .phase_sync_strobe_i(n533),
    .phase_set_strobe_i(n534),
    .phase_value_i(n535),
    .wave_o(\gen_channels_n7_channel_inst.wave_o ));
  /* ../../vhdl/src/synthesizer.vhd:25:55  */
  assign n532 = phase_increment_i[63:32]; // extract
  /* ../../vhdl/src/synthesizer.vhd:26:59  */
  assign n533 = phase_sync_strobe_i[6]; // extract
  /* ../../vhdl/src/synthesizer.vhd:27:57  */
  assign n534 = phase_set_strobe_i[6]; // extract
  /* ../../vhdl/src/synthesizer.vhd:28:47  */
  assign n535 = phase_value_i[63:32]; // extract
  /* ../../vhdl/src/synthesizer.vhd:21:9  */
  channel gen_channels_n8_channel_inst (
    .clock_i(clock_i),
    .reset_i(reset_i),
    .phase_increment_i(n537),
    .phase_sync_strobe_i(n538),
    .phase_set_strobe_i(n539),
    .phase_value_i(n540),
    .wave_o(\gen_channels_n8_channel_inst.wave_o ));
  /* ../../vhdl/src/synthesizer.vhd:25:55  */
  assign n537 = phase_increment_i[31:0]; // extract
  /* ../../vhdl/src/synthesizer.vhd:26:59  */
  assign n538 = phase_sync_strobe_i[7]; // extract
  /* ../../vhdl/src/synthesizer.vhd:27:57  */
  assign n539 = phase_set_strobe_i[7]; // extract
  /* ../../vhdl/src/synthesizer.vhd:28:47  */
  assign n540 = phase_value_i[31:0]; // extract
  assign n542 = {\gen_channels_n8_channel_inst.wave_o , \gen_channels_n7_channel_inst.wave_o , \gen_channels_n6_channel_inst.wave_o , \gen_channels_n5_channel_inst.wave_o , \gen_channels_n4_channel_inst.wave_o , \gen_channels_n3_channel_inst.wave_o , \gen_channels_n2_channel_inst.wave_o , \gen_channels_n1_channel_inst.wave_o };
endmodule

module uart_decoder
  (input  clock_i,
   input  reset_i,
   input  [7:0] rx_data_i,
   input  rx_valid_i,
   input  tx_busy_i,
   output [255:0] phase_increment_o,
   output [255:0] phase_value_o,
   output [7:0] phase_sync_strobe_o,
   output [7:0] phase_set_strobe_o,
   output [7:0] tx_data_o,
   output tx_valid_o);
  wire [7:0] rx_data_in_reg;
  wire rx_valid_in_reg;
  wire [2:0] rx_state_reg;
  wire [2:0] rx_state_next;
  wire [7:0] address_reg;
  wire [7:0] address_next;
  wire [7:0] instruction_reg;
  wire [7:0] instruction_next;
  wire [7:0] data1_reg;
  wire [7:0] data1_next;
  wire [7:0] data2_reg;
  wire [7:0] data2_next;
  wire [7:0] data3_reg;
  wire [7:0] data3_next;
  wire [7:0] data4_reg;
  wire [7:0] data4_next;
  wire [255:0] phase_inc_regs;
  wire [255:0] phase_inc_next;
  wire [255:0] phase_val_regs;
  wire [255:0] phase_val_next;
  wire [7:0] sync_strobe_reg;
  wire [7:0] sync_strobe_next;
  wire [7:0] set_strobe_reg;
  wire [7:0] set_strobe_next;
  wire [2:0] tx_state_reg;
  wire [2:0] tx_state_next;
  wire [7:0] tx_data_reg;
  wire [7:0] tx_data_next;
  wire tx_valid_reg;
  wire tx_valid_next;
  wire tx_busy_prev_reg;
  wire tx_start_reg;
  wire tx_start_next;
  wire n83;
  wire n84;
  wire n87;
  wire n90;
  wire [2:0] n92;
  wire n94;
  wire n96;
  wire n98;
  wire n100;
  wire n102;
  wire n104;
  wire n106;
  wire n108;
  wire n110;
  wire n112;
  wire n113;
  wire n115;
  wire [31:0] n117;
  wire n119;
  wire [31:0] n120;
  wire n122;
  wire n123;
  wire [31:0] n124;
  wire [31:0] n126;
  wire [2:0] n127;
  wire [15:0] n128;
  wire [23:0] n129;
  wire [31:0] n130;
  wire [2:0] n132;
  wire n136;
  localparam [7:0] n138 = 8'b00000000;
  wire n142;
  wire [2:0] n144;
  localparam [7:0] n148 = 8'b00000000;
  wire n152;
  wire [2:0] n153;
  reg [255:0] n154;
  reg [255:0] n155;
  reg [7:0] n157;
  reg [7:0] n159;
  wire [255:0] n160;
  wire [255:0] n161;
  wire [7:0] n163;
  wire [7:0] n165;
  wire n168;
  wire n169;
  wire [7:0] n171;
  wire [7:0] n173;
  wire n174;
  wire n179;
  wire [7:0] n180;
  reg [2:0] n189;
  reg [7:0] n190;
  reg [7:0] n191;
  reg [7:0] n192;
  reg [7:0] n193;
  reg [7:0] n194;
  reg [7:0] n195;
  reg [255:0] n196;
  reg [255:0] n197;
  reg [7:0] n199;
  reg [7:0] n201;
  reg n202;
  wire [2:0] n206;
  wire [7:0] n207;
  wire [7:0] n208;
  wire [7:0] n209;
  wire [7:0] n210;
  wire [7:0] n211;
  wire [7:0] n212;
  wire [255:0] n213;
  wire [255:0] n214;
  wire [7:0] n216;
  wire [7:0] n219;
  wire n221;
  wire n225;
  wire n226;
  wire [2:0] n228;
  wire [7:0] n229;
  wire n232;
  wire n234;
  wire n236;
  wire [2:0] n238;
  wire [7:0] n239;
  wire n242;
  wire n244;
  wire [2:0] n246;
  wire [7:0] n247;
  wire n250;
  wire n252;
  wire [2:0] n254;
  wire [7:0] n255;
  wire n258;
  wire n260;
  wire [2:0] n262;
  wire [7:0] n263;
  wire n266;
  wire n268;
  wire [2:0] n270;
  wire [7:0] n271;
  wire n274;
  wire n276;
  wire [5:0] n277;
  reg [2:0] n279;
  reg [7:0] n280;
  reg n282;
  reg n284;
  reg [7:0] n343;
  reg n344;
  reg [2:0] n345;
  reg [7:0] n346;
  reg [7:0] n347;
  reg [7:0] n348;
  reg [7:0] n349;
  reg [7:0] n350;
  reg [7:0] n351;
  reg [255:0] n352;
  reg [255:0] n353;
  reg [7:0] n354;
  reg [7:0] n355;
  reg [2:0] n356;
  reg [7:0] n357;
  reg n358;
  reg n359;
  reg n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire [31:0] n379;
  wire [31:0] n380;
  wire [31:0] n381;
  wire [31:0] n382;
  wire [31:0] n383;
  wire [31:0] n384;
  wire [31:0] n385;
  wire [31:0] n386;
  wire [31:0] n387;
  wire [31:0] n388;
  wire [31:0] n389;
  wire [31:0] n390;
  wire [31:0] n391;
  wire [31:0] n392;
  wire [31:0] n393;
  wire [31:0] n394;
  wire [255:0] n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire [7:0] n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire [31:0] n449;
  wire [31:0] n450;
  wire [31:0] n451;
  wire [31:0] n452;
  wire [31:0] n453;
  wire [31:0] n454;
  wire [31:0] n455;
  wire [31:0] n456;
  wire [31:0] n457;
  wire [31:0] n458;
  wire [31:0] n459;
  wire [31:0] n460;
  wire [31:0] n461;
  wire [31:0] n462;
  wire [31:0] n463;
  wire [31:0] n464;
  wire [255:0] n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire [7:0] n500;
  assign phase_increment_o = phase_inc_regs; //(module output)
  assign phase_value_o = phase_val_regs; //(module output)
  assign phase_sync_strobe_o = sync_strobe_reg; //(module output)
  assign phase_set_strobe_o = set_strobe_reg; //(module output)
  assign tx_data_o = tx_data_reg; //(module output)
  assign tx_valid_o = tx_valid_reg; //(module output)
  /* ../../vhdl/src/UART_DECODER.vhd:24:10  */
  assign rx_data_in_reg = n343; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:25:10  */
  assign rx_valid_in_reg = n344; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:28:10  */
  assign rx_state_reg = n345; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:29:10  */
  assign rx_state_next = n206; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:31:10  */
  assign address_reg = n346; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:32:10  */
  assign address_next = n207; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:33:10  */
  assign instruction_reg = n347; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:34:10  */
  assign instruction_next = n208; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:35:10  */
  assign data1_reg = n348; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:36:10  */
  assign data1_next = n209; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:37:10  */
  assign data2_reg = n349; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:38:10  */
  assign data2_next = n210; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:39:10  */
  assign data3_reg = n350; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:40:10  */
  assign data3_next = n211; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:41:10  */
  assign data4_reg = n351; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:42:10  */
  assign data4_next = n212; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:44:10  */
  assign phase_inc_regs = n352; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:45:10  */
  assign phase_inc_next = n213; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:46:10  */
  assign phase_val_regs = n353; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:47:10  */
  assign phase_val_next = n214; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:49:10  */
  assign sync_strobe_reg = n354; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:50:10  */
  assign sync_strobe_next = n216; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:51:10  */
  assign set_strobe_reg = n355; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:52:10  */
  assign set_strobe_next = n219; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:55:10  */
  assign tx_state_reg = n356; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:56:10  */
  assign tx_state_next = n279; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:57:10  */
  assign tx_data_reg = n357; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:58:10  */
  assign tx_data_next = n280; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:59:10  */
  assign tx_valid_reg = n358; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:60:10  */
  assign tx_valid_next = n282; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:61:10  */
  assign tx_busy_prev_reg = n359; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:62:10  */
  assign tx_start_reg = n360; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:63:10  */
  assign tx_start_next = n284; // (signal)
  /* ../../vhdl/src/UART_DECODER.vhd:95:48  */
  assign n83 = ~tx_busy_i;
  /* ../../vhdl/src/UART_DECODER.vhd:95:33  */
  assign n84 = n83 & tx_busy_prev_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:95:5  */
  assign n87 = n84 ? 1'b1 : 1'b0;
  /* ../../vhdl/src/UART_DECODER.vhd:102:29  */
  assign n90 = rx_data_in_reg == 8'b10101010;
  /* ../../vhdl/src/UART_DECODER.vhd:102:11  */
  assign n92 = n90 ? 3'b001 : rx_state_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:101:9  */
  assign n94 = rx_state_reg == 3'b000;
  /* ../../vhdl/src/UART_DECODER.vhd:105:9  */
  assign n96 = rx_state_reg == 3'b001;
  /* ../../vhdl/src/UART_DECODER.vhd:108:9  */
  assign n98 = rx_state_reg == 3'b010;
  /* ../../vhdl/src/UART_DECODER.vhd:111:9  */
  assign n100 = rx_state_reg == 3'b011;
  /* ../../vhdl/src/UART_DECODER.vhd:114:9  */
  assign n102 = rx_state_reg == 3'b100;
  /* ../../vhdl/src/UART_DECODER.vhd:117:9  */
  assign n104 = rx_state_reg == 3'b101;
  /* ../../vhdl/src/UART_DECODER.vhd:120:9  */
  assign n106 = rx_state_reg == 3'b110;
  /* ../../vhdl/src/UART_DECODER.vhd:124:29  */
  assign n108 = rx_data_in_reg == 8'b01010101;
  /* ../../vhdl/src/UART_DECODER.vhd:126:29  */
  assign n110 = address_reg == 8'b00000000;
  /* ../../vhdl/src/UART_DECODER.vhd:126:57  */
  assign n112 = instruction_reg == 8'b00000000;
  /* ../../vhdl/src/UART_DECODER.vhd:126:37  */
  assign n113 = n112 & n110;
  /* ../../vhdl/src/UART_DECODER.vhd:124:11  */
  assign n115 = n174 ? 1'b1 : tx_start_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:132:27  */
  assign n117 = {24'b0, address_reg};  //  uext
  /* ../../vhdl/src/UART_DECODER.vhd:132:27  */
  assign n119 = $signed(n117) >= $signed(32'b00000000000000000000000000000001);
  /* ../../vhdl/src/UART_DECODER.vhd:132:47  */
  assign n120 = {24'b0, address_reg};  //  uext
  /* ../../vhdl/src/UART_DECODER.vhd:132:47  */
  assign n122 = $signed(n120) <= $signed(32'b00000000000000000000000000001000);
  /* ../../vhdl/src/UART_DECODER.vhd:132:33  */
  assign n123 = n122 & n119;
  /* ../../vhdl/src/UART_DECODER.vhd:133:41  */
  assign n124 = {24'b0, address_reg};  //  uext
  /* ../../vhdl/src/UART_DECODER.vhd:133:41  */
  assign n126 = n124 - 32'b00000000000000000000000000000001;
  /* ../../vhdl/src/UART_DECODER.vhd:133:17  */
  assign n127 = n126[2:0];  // trunc
  /* ../../vhdl/src/UART_DECODER.vhd:134:53  */
  assign n128 = {data1_reg, data2_reg};
  /* ../../vhdl/src/UART_DECODER.vhd:134:65  */
  assign n129 = {n128, data3_reg};
  /* ../../vhdl/src/UART_DECODER.vhd:134:77  */
  assign n130 = {n129, data4_reg};
  /* ../../vhdl/src/UART_DECODER.vhd:138:40  */
  assign n132 = 3'b111 - n127;
  /* ../../vhdl/src/UART_DECODER.vhd:137:21  */
  assign n136 = instruction_reg == 8'b00000000;
  /* ../../vhdl/src/UART_DECODER.vhd:139:21  */
  assign n142 = instruction_reg == 8'b00000001;
  /* ../../vhdl/src/UART_DECODER.vhd:142:40  */
  assign n144 = 3'b111 - n127;
  /* ../../vhdl/src/UART_DECODER.vhd:141:21  */
  assign n152 = instruction_reg == 8'b00000010;
  assign n153 = {n152, n142, n136};
  /* ../../vhdl/src/UART_DECODER.vhd:136:17  */
  always @*
    case (n153)
      3'b100: n154 = phase_inc_regs;
      3'b010: n154 = phase_inc_regs;
      3'b001: n154 = n395;
      default: n154 = phase_inc_regs;
    endcase
  /* ../../vhdl/src/UART_DECODER.vhd:136:17  */
  always @*
    case (n153)
      3'b100: n155 = n465;
      3'b010: n155 = phase_val_regs;
      3'b001: n155 = phase_val_regs;
      default: n155 = phase_val_regs;
    endcase
  /* ../../vhdl/src/UART_DECODER.vhd:136:17  */
  always @*
    case (n153)
      3'b100: n157 = 8'b00000000;
      3'b010: n157 = n430;
      3'b001: n157 = 8'b00000000;
      default: n157 = 8'b00000000;
    endcase
  /* ../../vhdl/src/UART_DECODER.vhd:136:17  */
  always @*
    case (n153)
      3'b100: n159 = n500;
      3'b010: n159 = 8'b00000000;
      3'b001: n159 = 8'b00000000;
      default: n159 = 8'b00000000;
    endcase
  /* ../../vhdl/src/UART_DECODER.vhd:124:11  */
  assign n160 = n168 ? n154 : phase_inc_regs;
  /* ../../vhdl/src/UART_DECODER.vhd:124:11  */
  assign n161 = n169 ? n155 : phase_val_regs;
  /* ../../vhdl/src/UART_DECODER.vhd:132:14  */
  assign n163 = n123 ? n157 : 8'b00000000;
  /* ../../vhdl/src/UART_DECODER.vhd:132:14  */
  assign n165 = n123 ? n159 : 8'b00000000;
  /* ../../vhdl/src/UART_DECODER.vhd:124:11  */
  assign n168 = n123 & n108;
  /* ../../vhdl/src/UART_DECODER.vhd:124:11  */
  assign n169 = n123 & n108;
  /* ../../vhdl/src/UART_DECODER.vhd:124:11  */
  assign n171 = n108 ? n163 : 8'b00000000;
  /* ../../vhdl/src/UART_DECODER.vhd:124:11  */
  assign n173 = n108 ? n165 : 8'b00000000;
  /* ../../vhdl/src/UART_DECODER.vhd:124:11  */
  assign n174 = n113 & n108;
  /* ../../vhdl/src/UART_DECODER.vhd:123:9  */
  assign n179 = rx_state_reg == 3'b111;
  assign n180 = {n179, n106, n104, n102, n100, n98, n96, n94};
  /* ../../vhdl/src/UART_DECODER.vhd:100:7  */
  always @*
    case (n180)
      8'b10000000: n189 = 3'b000;
      8'b01000000: n189 = 3'b111;
      8'b00100000: n189 = 3'b110;
      8'b00010000: n189 = 3'b101;
      8'b00001000: n189 = 3'b100;
      8'b00000100: n189 = 3'b011;
      8'b00000010: n189 = 3'b010;
      8'b00000001: n189 = n92;
      default: n189 = 3'b000;
    endcase
  /* ../../vhdl/src/UART_DECODER.vhd:100:7  */
  always @*
    case (n180)
      8'b10000000: n190 = address_reg;
      8'b01000000: n190 = address_reg;
      8'b00100000: n190 = address_reg;
      8'b00010000: n190 = address_reg;
      8'b00001000: n190 = address_reg;
      8'b00000100: n190 = address_reg;
      8'b00000010: n190 = rx_data_in_reg;
      8'b00000001: n190 = address_reg;
      default: n190 = address_reg;
    endcase
  /* ../../vhdl/src/UART_DECODER.vhd:100:7  */
  always @*
    case (n180)
      8'b10000000: n191 = instruction_reg;
      8'b01000000: n191 = instruction_reg;
      8'b00100000: n191 = instruction_reg;
      8'b00010000: n191 = instruction_reg;
      8'b00001000: n191 = instruction_reg;
      8'b00000100: n191 = rx_data_in_reg;
      8'b00000010: n191 = instruction_reg;
      8'b00000001: n191 = instruction_reg;
      default: n191 = instruction_reg;
    endcase
  /* ../../vhdl/src/UART_DECODER.vhd:100:7  */
  always @*
    case (n180)
      8'b10000000: n192 = data1_reg;
      8'b01000000: n192 = data1_reg;
      8'b00100000: n192 = data1_reg;
      8'b00010000: n192 = data1_reg;
      8'b00001000: n192 = rx_data_in_reg;
      8'b00000100: n192 = data1_reg;
      8'b00000010: n192 = data1_reg;
      8'b00000001: n192 = data1_reg;
      default: n192 = data1_reg;
    endcase
  /* ../../vhdl/src/UART_DECODER.vhd:100:7  */
  always @*
    case (n180)
      8'b10000000: n193 = data2_reg;
      8'b01000000: n193 = data2_reg;
      8'b00100000: n193 = data2_reg;
      8'b00010000: n193 = rx_data_in_reg;
      8'b00001000: n193 = data2_reg;
      8'b00000100: n193 = data2_reg;
      8'b00000010: n193 = data2_reg;
      8'b00000001: n193 = data2_reg;
      default: n193 = data2_reg;
    endcase
  /* ../../vhdl/src/UART_DECODER.vhd:100:7  */
  always @*
    case (n180)
      8'b10000000: n194 = data3_reg;
      8'b01000000: n194 = data3_reg;
      8'b00100000: n194 = rx_data_in_reg;
      8'b00010000: n194 = data3_reg;
      8'b00001000: n194 = data3_reg;
      8'b00000100: n194 = data3_reg;
      8'b00000010: n194 = data3_reg;
      8'b00000001: n194 = data3_reg;
      default: n194 = data3_reg;
    endcase
  /* ../../vhdl/src/UART_DECODER.vhd:100:7  */
  always @*
    case (n180)
      8'b10000000: n195 = data4_reg;
      8'b01000000: n195 = rx_data_in_reg;
      8'b00100000: n195 = data4_reg;
      8'b00010000: n195 = data4_reg;
      8'b00001000: n195 = data4_reg;
      8'b00000100: n195 = data4_reg;
      8'b00000010: n195 = data4_reg;
      8'b00000001: n195 = data4_reg;
      default: n195 = data4_reg;
    endcase
  /* ../../vhdl/src/UART_DECODER.vhd:100:7  */
  always @*
    case (n180)
      8'b10000000: n196 = n160;
      8'b01000000: n196 = phase_inc_regs;
      8'b00100000: n196 = phase_inc_regs;
      8'b00010000: n196 = phase_inc_regs;
      8'b00001000: n196 = phase_inc_regs;
      8'b00000100: n196 = phase_inc_regs;
      8'b00000010: n196 = phase_inc_regs;
      8'b00000001: n196 = phase_inc_regs;
      default: n196 = phase_inc_regs;
    endcase
  /* ../../vhdl/src/UART_DECODER.vhd:100:7  */
  always @*
    case (n180)
      8'b10000000: n197 = n161;
      8'b01000000: n197 = phase_val_regs;
      8'b00100000: n197 = phase_val_regs;
      8'b00010000: n197 = phase_val_regs;
      8'b00001000: n197 = phase_val_regs;
      8'b00000100: n197 = phase_val_regs;
      8'b00000010: n197 = phase_val_regs;
      8'b00000001: n197 = phase_val_regs;
      default: n197 = phase_val_regs;
    endcase
  /* ../../vhdl/src/UART_DECODER.vhd:100:7  */
  always @*
    case (n180)
      8'b10000000: n199 = n171;
      8'b01000000: n199 = 8'b00000000;
      8'b00100000: n199 = 8'b00000000;
      8'b00010000: n199 = 8'b00000000;
      8'b00001000: n199 = 8'b00000000;
      8'b00000100: n199 = 8'b00000000;
      8'b00000010: n199 = 8'b00000000;
      8'b00000001: n199 = 8'b00000000;
      default: n199 = 8'b00000000;
    endcase
  /* ../../vhdl/src/UART_DECODER.vhd:100:7  */
  always @*
    case (n180)
      8'b10000000: n201 = n173;
      8'b01000000: n201 = 8'b00000000;
      8'b00100000: n201 = 8'b00000000;
      8'b00010000: n201 = 8'b00000000;
      8'b00001000: n201 = 8'b00000000;
      8'b00000100: n201 = 8'b00000000;
      8'b00000010: n201 = 8'b00000000;
      8'b00000001: n201 = 8'b00000000;
      default: n201 = 8'b00000000;
    endcase
  /* ../../vhdl/src/UART_DECODER.vhd:100:7  */
  always @*
    case (n180)
      8'b10000000: n202 = n115;
      8'b01000000: n202 = tx_start_reg;
      8'b00100000: n202 = tx_start_reg;
      8'b00010000: n202 = tx_start_reg;
      8'b00001000: n202 = tx_start_reg;
      8'b00000100: n202 = tx_start_reg;
      8'b00000010: n202 = tx_start_reg;
      8'b00000001: n202 = tx_start_reg;
      default: n202 = tx_start_reg;
    endcase
  /* ../../vhdl/src/UART_DECODER.vhd:99:5  */
  assign n206 = rx_valid_in_reg ? n189 : rx_state_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:99:5  */
  assign n207 = rx_valid_in_reg ? n190 : address_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:99:5  */
  assign n208 = rx_valid_in_reg ? n191 : instruction_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:99:5  */
  assign n209 = rx_valid_in_reg ? n192 : data1_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:99:5  */
  assign n210 = rx_valid_in_reg ? n193 : data2_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:99:5  */
  assign n211 = rx_valid_in_reg ? n194 : data3_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:99:5  */
  assign n212 = rx_valid_in_reg ? n195 : data4_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:99:5  */
  assign n213 = rx_valid_in_reg ? n196 : phase_inc_regs;
  /* ../../vhdl/src/UART_DECODER.vhd:99:5  */
  assign n214 = rx_valid_in_reg ? n197 : phase_val_regs;
  /* ../../vhdl/src/UART_DECODER.vhd:99:5  */
  assign n216 = rx_valid_in_reg ? n199 : 8'b00000000;
  /* ../../vhdl/src/UART_DECODER.vhd:99:5  */
  assign n219 = rx_valid_in_reg ? n201 : 8'b00000000;
  /* ../../vhdl/src/UART_DECODER.vhd:99:5  */
  assign n221 = rx_valid_in_reg ? n202 : tx_start_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:157:48  */
  assign n225 = ~tx_busy_i;
  /* ../../vhdl/src/UART_DECODER.vhd:157:33  */
  assign n226 = n225 & tx_start_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:157:9  */
  assign n228 = n226 ? 3'b001 : tx_state_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:157:9  */
  assign n229 = n226 ? address_reg : tx_data_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:157:9  */
  assign n232 = n226 ? 1'b1 : 1'b0;
  /* ../../vhdl/src/UART_DECODER.vhd:157:9  */
  assign n234 = n226 ? 1'b0 : n221;
  /* ../../vhdl/src/UART_DECODER.vhd:156:7  */
  assign n236 = tx_state_reg == 3'b000;
  /* ../../vhdl/src/UART_DECODER.vhd:164:9  */
  assign n238 = n87 ? 3'b010 : tx_state_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:164:9  */
  assign n239 = n87 ? instruction_reg : tx_data_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:164:9  */
  assign n242 = n87 ? 1'b1 : 1'b0;
  /* ../../vhdl/src/UART_DECODER.vhd:163:7  */
  assign n244 = tx_state_reg == 3'b001;
  /* ../../vhdl/src/UART_DECODER.vhd:170:9  */
  assign n246 = n87 ? 3'b011 : tx_state_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:170:9  */
  assign n247 = n87 ? data1_reg : tx_data_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:170:9  */
  assign n250 = n87 ? 1'b1 : 1'b0;
  /* ../../vhdl/src/UART_DECODER.vhd:169:7  */
  assign n252 = tx_state_reg == 3'b010;
  /* ../../vhdl/src/UART_DECODER.vhd:176:9  */
  assign n254 = n87 ? 3'b100 : tx_state_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:176:9  */
  assign n255 = n87 ? data2_reg : tx_data_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:176:9  */
  assign n258 = n87 ? 1'b1 : 1'b0;
  /* ../../vhdl/src/UART_DECODER.vhd:175:7  */
  assign n260 = tx_state_reg == 3'b011;
  /* ../../vhdl/src/UART_DECODER.vhd:182:9  */
  assign n262 = n87 ? 3'b101 : tx_state_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:182:9  */
  assign n263 = n87 ? data3_reg : tx_data_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:182:9  */
  assign n266 = n87 ? 1'b1 : 1'b0;
  /* ../../vhdl/src/UART_DECODER.vhd:181:7  */
  assign n268 = tx_state_reg == 3'b100;
  /* ../../vhdl/src/UART_DECODER.vhd:188:9  */
  assign n270 = n87 ? 3'b000 : tx_state_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:188:9  */
  assign n271 = n87 ? data4_reg : tx_data_reg;
  /* ../../vhdl/src/UART_DECODER.vhd:188:9  */
  assign n274 = n87 ? 1'b1 : 1'b0;
  /* ../../vhdl/src/UART_DECODER.vhd:187:7  */
  assign n276 = tx_state_reg == 3'b101;
  assign n277 = {n276, n268, n260, n252, n244, n236};
  /* ../../vhdl/src/UART_DECODER.vhd:155:5  */
  always @*
    case (n277)
      6'b100000: n279 = n270;
      6'b010000: n279 = n262;
      6'b001000: n279 = n254;
      6'b000100: n279 = n246;
      6'b000010: n279 = n238;
      6'b000001: n279 = n228;
      default: n279 = 3'b000;
    endcase
  /* ../../vhdl/src/UART_DECODER.vhd:155:5  */
  always @*
    case (n277)
      6'b100000: n280 = n271;
      6'b010000: n280 = n263;
      6'b001000: n280 = n255;
      6'b000100: n280 = n247;
      6'b000010: n280 = n239;
      6'b000001: n280 = n229;
      default: n280 = tx_data_reg;
    endcase
  /* ../../vhdl/src/UART_DECODER.vhd:155:5  */
  always @*
    case (n277)
      6'b100000: n282 = n274;
      6'b010000: n282 = n266;
      6'b001000: n282 = n258;
      6'b000100: n282 = n250;
      6'b000010: n282 = n242;
      6'b000001: n282 = n232;
      default: n282 = 1'b0;
    endcase
  /* ../../vhdl/src/UART_DECODER.vhd:155:5  */
  always @*
    case (n277)
      6'b100000: n284 = n221;
      6'b010000: n284 = n221;
      6'b001000: n284 = n221;
      6'b000100: n284 = n221;
      6'b000010: n284 = n221;
      6'b000001: n284 = n234;
      default: n284 = n221;
    endcase
  /* ../../vhdl/src/UART_DECODER.vhd:219:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n343 <= 8'b00000000;
    else
      n343 <= rx_data_i;
  /* ../../vhdl/src/UART_DECODER.vhd:219:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n344 <= 1'b0;
    else
      n344 <= rx_valid_i;
  /* ../../vhdl/src/UART_DECODER.vhd:219:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n345 <= 3'b000;
    else
      n345 <= rx_state_next;
  /* ../../vhdl/src/UART_DECODER.vhd:219:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n346 <= 8'b00000000;
    else
      n346 <= address_next;
  /* ../../vhdl/src/UART_DECODER.vhd:219:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n347 <= 8'b00000000;
    else
      n347 <= instruction_next;
  /* ../../vhdl/src/UART_DECODER.vhd:219:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n348 <= 8'b00000000;
    else
      n348 <= data1_next;
  /* ../../vhdl/src/UART_DECODER.vhd:219:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n349 <= 8'b00000000;
    else
      n349 <= data2_next;
  /* ../../vhdl/src/UART_DECODER.vhd:219:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n350 <= 8'b00000000;
    else
      n350 <= data3_next;
  /* ../../vhdl/src/UART_DECODER.vhd:219:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n351 <= 8'b00000000;
    else
      n351 <= data4_next;
  /* ../../vhdl/src/UART_DECODER.vhd:219:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n352 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n352 <= phase_inc_next;
  /* ../../vhdl/src/UART_DECODER.vhd:219:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n353 <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n353 <= phase_val_next;
  /* ../../vhdl/src/UART_DECODER.vhd:219:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n354 <= 8'b00000000;
    else
      n354 <= sync_strobe_next;
  /* ../../vhdl/src/UART_DECODER.vhd:219:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n355 <= 8'b00000000;
    else
      n355 <= set_strobe_next;
  /* ../../vhdl/src/UART_DECODER.vhd:219:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n356 <= 3'b000;
    else
      n356 <= tx_state_next;
  /* ../../vhdl/src/UART_DECODER.vhd:219:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n357 <= 8'b00000000;
    else
      n357 <= tx_data_next;
  /* ../../vhdl/src/UART_DECODER.vhd:219:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n358 <= 1'b0;
    else
      n358 <= tx_valid_next;
  /* ../../vhdl/src/UART_DECODER.vhd:219:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n359 <= 1'b0;
    else
      n359 <= tx_busy_i;
  /* ../../vhdl/src/UART_DECODER.vhd:219:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n360 <= 1'b0;
    else
      n360 <= tx_start_next;
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n361 = n132[2]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n362 = ~n361;
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n363 = n132[1]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n364 = ~n363;
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n365 = n362 & n364;
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n366 = n362 & n363;
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n367 = n361 & n364;
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n368 = n361 & n363;
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n369 = n132[0]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n370 = ~n369;
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n371 = n365 & n370;
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n372 = n365 & n369;
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n373 = n366 & n370;
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n374 = n366 & n369;
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n375 = n367 & n370;
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n376 = n367 & n369;
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n377 = n368 & n370;
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n378 = n368 & n369;
  /* ../../vhdl/src/UART_DECODER.vhd:200:5  */
  assign n379 = phase_inc_regs[31:0]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n380 = n371 ? n130 : n379;
  /* ../../vhdl/src/UART_DECODER.vhd:200:5  */
  assign n381 = phase_inc_regs[63:32]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n382 = n372 ? n130 : n381;
  /* ../../vhdl/src/UART_DECODER.vhd:200:5  */
  assign n383 = phase_inc_regs[95:64]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n384 = n373 ? n130 : n383;
  assign n385 = phase_inc_regs[127:96]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n386 = n374 ? n130 : n385;
  assign n387 = phase_inc_regs[159:128]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n388 = n375 ? n130 : n387;
  /* ../../vhdl/src/UART_DECODER.vhd:99:5  */
  assign n389 = phase_inc_regs[191:160]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n390 = n376 ? n130 : n389;
  /* ../../vhdl/src/UART_DECODER.vhd:99:5  */
  assign n391 = phase_inc_regs[223:192]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n392 = n377 ? n130 : n391;
  assign n393 = phase_inc_regs[255:224]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:138:25  */
  assign n394 = n378 ? n130 : n393;
  /* ../../vhdl/src/UART_DECODER.vhd:100:7  */
  assign n395 = {n394, n392, n390, n388, n386, n384, n382, n380};
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n396 = n127[2]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n397 = ~n396;
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n398 = n127[1]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n399 = ~n398;
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n400 = n397 & n399;
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n401 = n397 & n398;
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n402 = n396 & n399;
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n403 = n396 & n398;
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n404 = n127[0]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n405 = ~n404;
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n406 = n400 & n405;
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n407 = n400 & n404;
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n408 = n401 & n405;
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n409 = n401 & n404;
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n410 = n402 & n405;
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n411 = n402 & n404;
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n412 = n403 & n405;
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n413 = n403 & n404;
  assign n414 = n138[0]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n415 = n406 ? 1'b1 : n414;
  assign n416 = n138[1]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n417 = n407 ? 1'b1 : n416;
  assign n418 = n138[2]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n419 = n408 ? 1'b1 : n418;
  assign n420 = n138[3]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n421 = n409 ? 1'b1 : n420;
  assign n422 = n138[4]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n423 = n410 ? 1'b1 : n422;
  assign n424 = n138[5]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n425 = n411 ? 1'b1 : n424;
  assign n426 = n138[6]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n427 = n412 ? 1'b1 : n426;
  assign n428 = n138[7]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:140:25  */
  assign n429 = n413 ? 1'b1 : n428;
  assign n430 = {n429, n427, n425, n423, n421, n419, n417, n415};
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n431 = n144[2]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n432 = ~n431;
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n433 = n144[1]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n434 = ~n433;
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n435 = n432 & n434;
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n436 = n432 & n433;
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n437 = n431 & n434;
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n438 = n431 & n433;
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n439 = n144[0]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n440 = ~n439;
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n441 = n435 & n440;
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n442 = n435 & n439;
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n443 = n436 & n440;
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n444 = n436 & n439;
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n445 = n437 & n440;
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n446 = n437 & n439;
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n447 = n438 & n440;
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n448 = n438 & n439;
  assign n449 = phase_val_regs[31:0]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n450 = n441 ? n130 : n449;
  assign n451 = phase_val_regs[63:32]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n452 = n442 ? n130 : n451;
  assign n453 = phase_val_regs[95:64]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n454 = n443 ? n130 : n453;
  assign n455 = phase_val_regs[127:96]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n456 = n444 ? n130 : n455;
  assign n457 = phase_val_regs[159:128]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n458 = n445 ? n130 : n457;
  assign n459 = phase_val_regs[191:160]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n460 = n446 ? n130 : n459;
  assign n461 = phase_val_regs[223:192]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n462 = n447 ? n130 : n461;
  assign n463 = phase_val_regs[255:224]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:142:25  */
  assign n464 = n448 ? n130 : n463;
  assign n465 = {n464, n462, n460, n458, n456, n454, n452, n450};
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n466 = n127[2]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n467 = ~n466;
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n468 = n127[1]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n469 = ~n468;
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n470 = n467 & n469;
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n471 = n467 & n468;
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n472 = n466 & n469;
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n473 = n466 & n468;
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n474 = n127[0]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n475 = ~n474;
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n476 = n470 & n475;
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n477 = n470 & n474;
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n478 = n471 & n475;
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n479 = n471 & n474;
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n480 = n472 & n475;
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n481 = n472 & n474;
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n482 = n473 & n475;
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n483 = n473 & n474;
  assign n484 = n148[0]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n485 = n476 ? 1'b1 : n484;
  assign n486 = n148[1]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n487 = n477 ? 1'b1 : n486;
  assign n488 = n148[2]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n489 = n478 ? 1'b1 : n488;
  assign n490 = n148[3]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n491 = n479 ? 1'b1 : n490;
  assign n492 = n148[4]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n493 = n480 ? 1'b1 : n492;
  assign n494 = n148[5]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n495 = n481 ? 1'b1 : n494;
  assign n496 = n148[6]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n497 = n482 ? 1'b1 : n496;
  assign n498 = n148[7]; // extract
  /* ../../vhdl/src/UART_DECODER.vhd:143:25  */
  assign n499 = n483 ? 1'b1 : n498;
  assign n500 = {n499, n497, n495, n493, n491, n489, n487, n485};
endmodule

module uart_core
  (input  clock_i,
   input  reset_i,
   input  serial_rx_i,
   output serial_tx_o,
   output [7:0] rx_data_o,
   output rx_valid_o,
   input  [7:0] tx_data_i,
   input  tx_valid_i,
   output tx_busy_o);
  wire rx_valid_sig;
  wire [7:0] rx_byte_sig;
  wire tx_data_valid_reg;
  wire tx_data_valid_next;
  wire [7:0] tx_byte_reg;
  wire [7:0] tx_byte_next;
  wire tx_done_sig;
  wire tx_state_reg;
  wire tx_state_next;
  wire tx_busy_reg;
  wire tx_busy_next;
  wire \uart_tx_inst.tx_active_o ;
  wire \uart_tx_inst.serial_o ;
  wire n25;
  wire [7:0] n26;
  wire n28;
  wire n31;
  wire n34;
  wire n37;
  wire n39;
  wire [1:0] n40;
  reg n43;
  reg [7:0] n46;
  reg n48;
  reg n51;
  reg n68;
  reg [7:0] n69;
  reg n70;
  reg n71;
  assign serial_tx_o = \uart_tx_inst.serial_o ; //(module output)
  assign rx_data_o = rx_byte_sig; //(module output)
  assign rx_valid_o = rx_valid_sig; //(module output)
  assign tx_busy_o = tx_busy_reg; //(module output)
  /* ../../vhdl/src/UART_CORE.vhd:24:10  */
  assign tx_data_valid_reg = n68; // (signal)
  /* ../../vhdl/src/UART_CORE.vhd:25:10  */
  assign tx_data_valid_next = n43; // (signal)
  /* ../../vhdl/src/UART_CORE.vhd:26:10  */
  assign tx_byte_reg = n69; // (signal)
  /* ../../vhdl/src/UART_CORE.vhd:27:10  */
  assign tx_byte_next = n46; // (signal)
  /* ../../vhdl/src/UART_CORE.vhd:30:10  */
  assign tx_state_reg = n70; // (signal)
  /* ../../vhdl/src/UART_CORE.vhd:31:10  */
  assign tx_state_next = n48; // (signal)
  /* ../../vhdl/src/UART_CORE.vhd:32:10  */
  assign tx_busy_reg = n71; // (signal)
  /* ../../vhdl/src/UART_CORE.vhd:33:10  */
  assign tx_busy_next = n51; // (signal)
  /* ../../vhdl/src/UART_CORE.vhd:37:3  */
  uart_rx uart_rx_inst (
    .clock_i(clock_i),
    .reset_i(reset_i),
    .serial_i(serial_rx_i),
    .data_valid_o(rx_valid_sig),
    .rx_byte_o(rx_byte_sig));
  /* ../../vhdl/src/UART_CORE.vhd:46:3  */
  uart_tx uart_tx_inst (
    .clock_i(clock_i),
    .reset_i(reset_i),
    .tx_data_valid_i(tx_data_valid_reg),
    .tx_data_i(tx_byte_reg),
    .tx_active_o(),
    .serial_o(\uart_tx_inst.serial_o ),
    .tx_done_o(tx_done_sig));
  /* ../../vhdl/src/UART_CORE.vhd:77:9  */
  assign n25 = tx_valid_i ? 1'b1 : 1'b0;
  /* ../../vhdl/src/UART_CORE.vhd:77:9  */
  assign n26 = tx_valid_i ? tx_data_i : tx_byte_reg;
  /* ../../vhdl/src/UART_CORE.vhd:77:9  */
  assign n28 = tx_valid_i ? 1'b1 : tx_state_reg;
  /* ../../vhdl/src/UART_CORE.vhd:77:9  */
  assign n31 = tx_valid_i ? 1'b1 : 1'b0;
  /* ../../vhdl/src/UART_CORE.vhd:74:7  */
  assign n34 = tx_state_reg == 1'b0;
  /* ../../vhdl/src/UART_CORE.vhd:88:9  */
  assign n37 = tx_done_sig ? 1'b0 : 1'b1;
  /* ../../vhdl/src/UART_CORE.vhd:84:7  */
  assign n39 = tx_state_reg == 1'b1;
  assign n40 = {n39, n34};
  /* ../../vhdl/src/UART_CORE.vhd:72:5  */
  always @*
    case (n40)
      2'b10: n43 = 1'b0;
      2'b01: n43 = n25;
      default: n43 = 1'b0;
    endcase
  /* ../../vhdl/src/UART_CORE.vhd:72:5  */
  always @*
    case (n40)
      2'b10: n46 = tx_byte_reg;
      2'b01: n46 = n26;
      default: n46 = 8'b00000000;
    endcase
  /* ../../vhdl/src/UART_CORE.vhd:72:5  */
  always @*
    case (n40)
      2'b10: n48 = n37;
      2'b01: n48 = n28;
      default: n48 = 1'b0;
    endcase
  /* ../../vhdl/src/UART_CORE.vhd:72:5  */
  always @*
    case (n40)
      2'b10: n51 = 1'b1;
      2'b01: n51 = n31;
      default: n51 = 1'b1;
    endcase
  /* ../../vhdl/src/UART_CORE.vhd:110:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n68 <= 1'b0;
    else
      n68 <= tx_data_valid_next;
  /* ../../vhdl/src/UART_CORE.vhd:110:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n69 <= 8'b00000000;
    else
      n69 <= tx_byte_next;
  /* ../../vhdl/src/UART_CORE.vhd:110:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n70 <= 1'b0;
    else
      n70 <= tx_state_next;
  /* ../../vhdl/src/UART_CORE.vhd:110:5  */
  always @(posedge clock_i or posedge reset_i)
    if (reset_i)
      n71 <= 1'b0;
    else
      n71 <= tx_busy_next;
endmodule

module octawave
  (input  clock_i,
   input  reset_n_i,
   input  uart_rx,
   output uart_tx,
   output [7:0] channel_o);
  wire reset;
  wire [7:0] rx_data;
  wire rx_valid;
  wire [7:0] tx_data;
  wire tx_valid;
  wire tx_busy;
  wire [255:0] phase_increment;
  wire [255:0] phase_value;
  wire [7:0] phase_sync_strobe;
  wire [7:0] phase_set_strobe;
  wire [7:0] waves;
  wire n2;
  wire \uart_core_inst.serial_tx_o ;
  assign uart_tx = \uart_core_inst.serial_tx_o ; //(module output)
  assign channel_o = waves; //(module output)
  /* ../../vhdl/src/octawave.vhd:17:10  */
  assign reset = n2; // (signal)
  /* ../../vhdl/src/octawave.vhd:32:12  */
  assign n2 = ~reset_n_i;
  /* ../../vhdl/src/octawave.vhd:34:3  */
  uart_core uart_core_inst (
    .clock_i(clock_i),
    .reset_i(reset),
    .serial_rx_i(uart_rx),
    .tx_data_i(tx_data),
    .tx_valid_i(tx_valid),
    .serial_tx_o(\uart_core_inst.serial_tx_o ),
    .rx_data_o(rx_data),
    .rx_valid_o(rx_valid),
    .tx_busy_o(tx_busy));
  /* ../../vhdl/src/octawave.vhd:47:3  */
  uart_decoder uart_decoder_inst (
    .clock_i(clock_i),
    .reset_i(reset),
    .rx_data_i(rx_data),
    .rx_valid_i(rx_valid),
    .tx_busy_i(tx_busy),
    .phase_increment_o(phase_increment),
    .phase_value_o(phase_value),
    .phase_sync_strobe_o(phase_sync_strobe),
    .phase_set_strobe_o(phase_set_strobe),
    .tx_data_o(tx_data),
    .tx_valid_o(tx_valid));
  /* ../../vhdl/src/octawave.vhd:62:3  */
  synthesizer synthesizer_inst (
    .clock_i(clock_i),
    .reset_i(reset),
    .phase_increment_i(phase_increment),
    .phase_value_i(phase_value),
    .phase_sync_strobe_i(phase_sync_strobe),
    .phase_set_strobe_i(phase_set_strobe),
    .waves_o(waves));
endmodule

